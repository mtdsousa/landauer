//Written by the Majority Logic Package Thu Jul  2 16:59:23 2015
module top (
            A_0, A_1, A_2, A_3, A_4, A_5, A_6, A_7, A_8, A_9, A_10, A_11, A_12, A_13, A_14, A_15, A_16, A_17, A_18, A_19, A_20, A_21, A_22, A_23, A_24, A_25, A_26, A_27, A_28, A_29, A_30, A_31, A_32, A_33, A_34, A_35, A_36, A_37, A_38, A_39, A_40, A_41, A_42, A_43, A_44, A_45, A_46, A_47, A_48, A_49, A_50, A_51, A_52, A_53, A_54, A_55, A_56, A_57, A_58, A_59, A_60, A_61, A_62, A_63, A_64, A_65, A_66, A_67, A_68, A_69, A_70, A_71, A_72, A_73, A_74, A_75, A_76, A_77, A_78, A_79, A_80, A_81, A_82, A_83, A_84, A_85, A_86, A_87, A_88, A_89, A_90, A_91, A_92, A_93, A_94, A_95, A_96, A_97, A_98, A_99, A_100, A_101, A_102, A_103, A_104, A_105, A_106, A_107, A_108, A_109, A_110, A_111, A_112, A_113, A_114, A_115, A_116, A_117, A_118, A_119, A_120, A_121, A_122, A_123, A_124, A_125, A_126, A_127, A_128, A_129, A_130, A_131, A_132, A_133, A_134, A_135, A_136, A_137, A_138, A_139, A_140, A_141, A_142, A_143, A_144, A_145, A_146, A_147, A_148, A_149, A_150, A_151, A_152, A_153, A_154, A_155, A_156, A_157, A_158, A_159, A_160, A_161, A_162, A_163, A_164, A_165, A_166, A_167, A_168, A_169, A_170, A_171, A_172, A_173, A_174, A_175, A_176, A_177, A_178, A_179, A_180, A_181, A_182, A_183, A_184, A_185, A_186, A_187, A_188, A_189, A_190, A_191, A_192, A_193, A_194, A_195, A_196, A_197, A_198, A_199, A_200, A_201, A_202, A_203, A_204, A_205, A_206, A_207, A_208, A_209, A_210, A_211, A_212, A_213, A_214, A_215, A_216, A_217, A_218, A_219, A_220, A_221, A_222, A_223, A_224, A_225, A_226, A_227, A_228, A_229, A_230, A_231, A_232, A_233, A_234, A_235, A_236, A_237, A_238, A_239, A_240, A_241, A_242, A_243, A_244, A_245, A_246, A_247, A_248, A_249, A_250, A_251, A_252, A_253, A_254, A_255, A_256, A_257, A_258, A_259, A_260, A_261, A_262, A_263, A_264, A_265, A_266, A_267, A_268, A_269, A_270, A_271, A_272, A_273, A_274, A_275, A_276, A_277, A_278, A_279, A_280, A_281, A_282, A_283, A_284, A_285, A_286, A_287, A_288, A_289, A_290, A_291, A_292, A_293, A_294, A_295, A_296, A_297, A_298, A_299, A_300, A_301, A_302, A_303, A_304, A_305, A_306, A_307, A_308, A_309, A_310, A_311, A_312, A_313, A_314, A_315, A_316, A_317, A_318, A_319, A_320, A_321, A_322, A_323, A_324, A_325, A_326, A_327, A_328, A_329, A_330, A_331, A_332, A_333, A_334, A_335, A_336, A_337, A_338, A_339, A_340, A_341, A_342, A_343, A_344, A_345, A_346, A_347, A_348, A_349, A_350, A_351, A_352, A_353, A_354, A_355, A_356, A_357, A_358, A_359, A_360, A_361, A_362, A_363, A_364, A_365, A_366, A_367, A_368, A_369, A_370, A_371, A_372, A_373, A_374, A_375, A_376, A_377, A_378, A_379, A_380, A_381, A_382, A_383, A_384, A_385, A_386, A_387, A_388, A_389, A_390, A_391, A_392, A_393, A_394, A_395, A_396, A_397, A_398, A_399, A_400, A_401, A_402, A_403, A_404, A_405, A_406, A_407, A_408, A_409, A_410, A_411, A_412, A_413, A_414, A_415, A_416, A_417, A_418, A_419, A_420, A_421, A_422, A_423, A_424, A_425, A_426, A_427, A_428, A_429, A_430, A_431, A_432, A_433, A_434, A_435, A_436, A_437, A_438, A_439, A_440, A_441, A_442, A_443, A_444, A_445, A_446, A_447, A_448, A_449, A_450, A_451, A_452, A_453, A_454, A_455, A_456, A_457, A_458, A_459, A_460, A_461, A_462, A_463, A_464, A_465, A_466, A_467, A_468, A_469, A_470, A_471, A_472, A_473, A_474, A_475, A_476, A_477, A_478, A_479, A_480, A_481, A_482, A_483, A_484, A_485, A_486, A_487, A_488, A_489, A_490, A_491, A_492, A_493, A_494, A_495, A_496, A_497, A_498, A_499, A_500, A_501, A_502, A_503, A_504, A_505, A_506, A_507, A_508, A_509, A_510, A_511, A_512, A_513, A_514, A_515, A_516, A_517, A_518, A_519, A_520, A_521, A_522, A_523, A_524, A_525, A_526, A_527, A_528, A_529, A_530, A_531, A_532, A_533, A_534, A_535, A_536, A_537, A_538, A_539, A_540, A_541, A_542, A_543, A_544, A_545, A_546, A_547, A_548, A_549, A_550, A_551, A_552, A_553, A_554, A_555, A_556, A_557, A_558, A_559, A_560, A_561, A_562, A_563, A_564, A_565, A_566, A_567, A_568, A_569, A_570, A_571, A_572, A_573, A_574, A_575, A_576, A_577, A_578, A_579, A_580, A_581, A_582, A_583, A_584, A_585, A_586, A_587, A_588, A_589, A_590, A_591, A_592, A_593, A_594, A_595, A_596, A_597, A_598, A_599, A_600, A_601, A_602, A_603, A_604, A_605, A_606, A_607, A_608, A_609, A_610, A_611, A_612, A_613, A_614, A_615, A_616, A_617, A_618, A_619, A_620, A_621, A_622, A_623, A_624, A_625, A_626, A_627, A_628, A_629, A_630, A_631, A_632, A_633, A_634, A_635, A_636, A_637, A_638, A_639, A_640, A_641, A_642, A_643, A_644, A_645, A_646, A_647, A_648, A_649, A_650, A_651, A_652, A_653, A_654, A_655, A_656, A_657, A_658, A_659, A_660, A_661, A_662, A_663, A_664, A_665, A_666, A_667, A_668, A_669, A_670, A_671, A_672, A_673, A_674, A_675, A_676, A_677, A_678, A_679, A_680, A_681, A_682, A_683, A_684, A_685, A_686, A_687, A_688, A_689, A_690, A_691, A_692, A_693, A_694, A_695, A_696, A_697, A_698, A_699, A_700, A_701, A_702, A_703, A_704, A_705, A_706, A_707, A_708, A_709, A_710, A_711, A_712, A_713, A_714, A_715, A_716, A_717, A_718, A_719, A_720, A_721, A_722, A_723, A_724, A_725, A_726, A_727, A_728, A_729, A_730, A_731, A_732, A_733, A_734, A_735, A_736, A_737, A_738, A_739, A_740, A_741, A_742, A_743, A_744, A_745, A_746, A_747, A_748, A_749, A_750, A_751, A_752, A_753, A_754, A_755, A_756, A_757, A_758, A_759, A_760, A_761, A_762, A_763, A_764, A_765, A_766, A_767, A_768, A_769, A_770, A_771, A_772, A_773, A_774, A_775, A_776, A_777, A_778, A_779, A_780, A_781, A_782, A_783, A_784, A_785, A_786, A_787, A_788, A_789, A_790, A_791, A_792, A_793, A_794, A_795, A_796, A_797, A_798, A_799, A_800, A_801, A_802, A_803, A_804, A_805, A_806, A_807, A_808, A_809, A_810, A_811, A_812, A_813, A_814, A_815, A_816, A_817, A_818, A_819, A_820, A_821, A_822, A_823, A_824, A_825, A_826, A_827, A_828, A_829, A_830, A_831, A_832, A_833, A_834, A_835, A_836, A_837, A_838, A_839, A_840, A_841, A_842, A_843, A_844, A_845, A_846, A_847, A_848, A_849, A_850, A_851, A_852, A_853, A_854, A_855, A_856, A_857, A_858, A_859, A_860, A_861, A_862, A_863, A_864, A_865, A_866, A_867, A_868, A_869, A_870, A_871, A_872, A_873, A_874, A_875, A_876, A_877, A_878, A_879, A_880, A_881, A_882, A_883, A_884, A_885, A_886, A_887, A_888, A_889, A_890, A_891, A_892, A_893, A_894, A_895, A_896, A_897, A_898, A_899, A_900, A_901, A_902, A_903, A_904, A_905, A_906, A_907, A_908, A_909, A_910, A_911, A_912, A_913, A_914, A_915, A_916, A_917, A_918, A_919, A_920, A_921, A_922, A_923, A_924, A_925, A_926, A_927, A_928, A_929, A_930, A_931, A_932, A_933, A_934, A_935, A_936, A_937, A_938, A_939, A_940, A_941, A_942, A_943, A_944, A_945, A_946, A_947, A_948, A_949, A_950, A_951, A_952, A_953, A_954, A_955, A_956, A_957, A_958, A_959, A_960, A_961, A_962, A_963, A_964, A_965, A_966, A_967, A_968, A_969, A_970, A_971, A_972, A_973, A_974, A_975, A_976, A_977, A_978, A_979, A_980, A_981, A_982, A_983, A_984, A_985, A_986, A_987, A_988, A_989, A_990, A_991, A_992, A_993, A_994, A_995, A_996, A_997, A_998, A_999, A_1000, 
            maj);
input A_0, A_1, A_2, A_3, A_4, A_5, A_6, A_7, A_8, A_9, A_10, A_11, A_12, A_13, A_14, A_15, A_16, A_17, A_18, A_19, A_20, A_21, A_22, A_23, A_24, A_25, A_26, A_27, A_28, A_29, A_30, A_31, A_32, A_33, A_34, A_35, A_36, A_37, A_38, A_39, A_40, A_41, A_42, A_43, A_44, A_45, A_46, A_47, A_48, A_49, A_50, A_51, A_52, A_53, A_54, A_55, A_56, A_57, A_58, A_59, A_60, A_61, A_62, A_63, A_64, A_65, A_66, A_67, A_68, A_69, A_70, A_71, A_72, A_73, A_74, A_75, A_76, A_77, A_78, A_79, A_80, A_81, A_82, A_83, A_84, A_85, A_86, A_87, A_88, A_89, A_90, A_91, A_92, A_93, A_94, A_95, A_96, A_97, A_98, A_99, A_100, A_101, A_102, A_103, A_104, A_105, A_106, A_107, A_108, A_109, A_110, A_111, A_112, A_113, A_114, A_115, A_116, A_117, A_118, A_119, A_120, A_121, A_122, A_123, A_124, A_125, A_126, A_127, A_128, A_129, A_130, A_131, A_132, A_133, A_134, A_135, A_136, A_137, A_138, A_139, A_140, A_141, A_142, A_143, A_144, A_145, A_146, A_147, A_148, A_149, A_150, A_151, A_152, A_153, A_154, A_155, A_156, A_157, A_158, A_159, A_160, A_161, A_162, A_163, A_164, A_165, A_166, A_167, A_168, A_169, A_170, A_171, A_172, A_173, A_174, A_175, A_176, A_177, A_178, A_179, A_180, A_181, A_182, A_183, A_184, A_185, A_186, A_187, A_188, A_189, A_190, A_191, A_192, A_193, A_194, A_195, A_196, A_197, A_198, A_199, A_200, A_201, A_202, A_203, A_204, A_205, A_206, A_207, A_208, A_209, A_210, A_211, A_212, A_213, A_214, A_215, A_216, A_217, A_218, A_219, A_220, A_221, A_222, A_223, A_224, A_225, A_226, A_227, A_228, A_229, A_230, A_231, A_232, A_233, A_234, A_235, A_236, A_237, A_238, A_239, A_240, A_241, A_242, A_243, A_244, A_245, A_246, A_247, A_248, A_249, A_250, A_251, A_252, A_253, A_254, A_255, A_256, A_257, A_258, A_259, A_260, A_261, A_262, A_263, A_264, A_265, A_266, A_267, A_268, A_269, A_270, A_271, A_272, A_273, A_274, A_275, A_276, A_277, A_278, A_279, A_280, A_281, A_282, A_283, A_284, A_285, A_286, A_287, A_288, A_289, A_290, A_291, A_292, A_293, A_294, A_295, A_296, A_297, A_298, A_299, A_300, A_301, A_302, A_303, A_304, A_305, A_306, A_307, A_308, A_309, A_310, A_311, A_312, A_313, A_314, A_315, A_316, A_317, A_318, A_319, A_320, A_321, A_322, A_323, A_324, A_325, A_326, A_327, A_328, A_329, A_330, A_331, A_332, A_333, A_334, A_335, A_336, A_337, A_338, A_339, A_340, A_341, A_342, A_343, A_344, A_345, A_346, A_347, A_348, A_349, A_350, A_351, A_352, A_353, A_354, A_355, A_356, A_357, A_358, A_359, A_360, A_361, A_362, A_363, A_364, A_365, A_366, A_367, A_368, A_369, A_370, A_371, A_372, A_373, A_374, A_375, A_376, A_377, A_378, A_379, A_380, A_381, A_382, A_383, A_384, A_385, A_386, A_387, A_388, A_389, A_390, A_391, A_392, A_393, A_394, A_395, A_396, A_397, A_398, A_399, A_400, A_401, A_402, A_403, A_404, A_405, A_406, A_407, A_408, A_409, A_410, A_411, A_412, A_413, A_414, A_415, A_416, A_417, A_418, A_419, A_420, A_421, A_422, A_423, A_424, A_425, A_426, A_427, A_428, A_429, A_430, A_431, A_432, A_433, A_434, A_435, A_436, A_437, A_438, A_439, A_440, A_441, A_442, A_443, A_444, A_445, A_446, A_447, A_448, A_449, A_450, A_451, A_452, A_453, A_454, A_455, A_456, A_457, A_458, A_459, A_460, A_461, A_462, A_463, A_464, A_465, A_466, A_467, A_468, A_469, A_470, A_471, A_472, A_473, A_474, A_475, A_476, A_477, A_478, A_479, A_480, A_481, A_482, A_483, A_484, A_485, A_486, A_487, A_488, A_489, A_490, A_491, A_492, A_493, A_494, A_495, A_496, A_497, A_498, A_499, A_500, A_501, A_502, A_503, A_504, A_505, A_506, A_507, A_508, A_509, A_510, A_511, A_512, A_513, A_514, A_515, A_516, A_517, A_518, A_519, A_520, A_521, A_522, A_523, A_524, A_525, A_526, A_527, A_528, A_529, A_530, A_531, A_532, A_533, A_534, A_535, A_536, A_537, A_538, A_539, A_540, A_541, A_542, A_543, A_544, A_545, A_546, A_547, A_548, A_549, A_550, A_551, A_552, A_553, A_554, A_555, A_556, A_557, A_558, A_559, A_560, A_561, A_562, A_563, A_564, A_565, A_566, A_567, A_568, A_569, A_570, A_571, A_572, A_573, A_574, A_575, A_576, A_577, A_578, A_579, A_580, A_581, A_582, A_583, A_584, A_585, A_586, A_587, A_588, A_589, A_590, A_591, A_592, A_593, A_594, A_595, A_596, A_597, A_598, A_599, A_600, A_601, A_602, A_603, A_604, A_605, A_606, A_607, A_608, A_609, A_610, A_611, A_612, A_613, A_614, A_615, A_616, A_617, A_618, A_619, A_620, A_621, A_622, A_623, A_624, A_625, A_626, A_627, A_628, A_629, A_630, A_631, A_632, A_633, A_634, A_635, A_636, A_637, A_638, A_639, A_640, A_641, A_642, A_643, A_644, A_645, A_646, A_647, A_648, A_649, A_650, A_651, A_652, A_653, A_654, A_655, A_656, A_657, A_658, A_659, A_660, A_661, A_662, A_663, A_664, A_665, A_666, A_667, A_668, A_669, A_670, A_671, A_672, A_673, A_674, A_675, A_676, A_677, A_678, A_679, A_680, A_681, A_682, A_683, A_684, A_685, A_686, A_687, A_688, A_689, A_690, A_691, A_692, A_693, A_694, A_695, A_696, A_697, A_698, A_699, A_700, A_701, A_702, A_703, A_704, A_705, A_706, A_707, A_708, A_709, A_710, A_711, A_712, A_713, A_714, A_715, A_716, A_717, A_718, A_719, A_720, A_721, A_722, A_723, A_724, A_725, A_726, A_727, A_728, A_729, A_730, A_731, A_732, A_733, A_734, A_735, A_736, A_737, A_738, A_739, A_740, A_741, A_742, A_743, A_744, A_745, A_746, A_747, A_748, A_749, A_750, A_751, A_752, A_753, A_754, A_755, A_756, A_757, A_758, A_759, A_760, A_761, A_762, A_763, A_764, A_765, A_766, A_767, A_768, A_769, A_770, A_771, A_772, A_773, A_774, A_775, A_776, A_777, A_778, A_779, A_780, A_781, A_782, A_783, A_784, A_785, A_786, A_787, A_788, A_789, A_790, A_791, A_792, A_793, A_794, A_795, A_796, A_797, A_798, A_799, A_800, A_801, A_802, A_803, A_804, A_805, A_806, A_807, A_808, A_809, A_810, A_811, A_812, A_813, A_814, A_815, A_816, A_817, A_818, A_819, A_820, A_821, A_822, A_823, A_824, A_825, A_826, A_827, A_828, A_829, A_830, A_831, A_832, A_833, A_834, A_835, A_836, A_837, A_838, A_839, A_840, A_841, A_842, A_843, A_844, A_845, A_846, A_847, A_848, A_849, A_850, A_851, A_852, A_853, A_854, A_855, A_856, A_857, A_858, A_859, A_860, A_861, A_862, A_863, A_864, A_865, A_866, A_867, A_868, A_869, A_870, A_871, A_872, A_873, A_874, A_875, A_876, A_877, A_878, A_879, A_880, A_881, A_882, A_883, A_884, A_885, A_886, A_887, A_888, A_889, A_890, A_891, A_892, A_893, A_894, A_895, A_896, A_897, A_898, A_899, A_900, A_901, A_902, A_903, A_904, A_905, A_906, A_907, A_908, A_909, A_910, A_911, A_912, A_913, A_914, A_915, A_916, A_917, A_918, A_919, A_920, A_921, A_922, A_923, A_924, A_925, A_926, A_927, A_928, A_929, A_930, A_931, A_932, A_933, A_934, A_935, A_936, A_937, A_938, A_939, A_940, A_941, A_942, A_943, A_944, A_945, A_946, A_947, A_948, A_949, A_950, A_951, A_952, A_953, A_954, A_955, A_956, A_957, A_958, A_959, A_960, A_961, A_962, A_963, A_964, A_965, A_966, A_967, A_968, A_969, A_970, A_971, A_972, A_973, A_974, A_975, A_976, A_977, A_978, A_979, A_980, A_981, A_982, A_983, A_984, A_985, A_986, A_987, A_988, A_989, A_990, A_991, A_992, A_993, A_994, A_995, A_996, A_997, A_998, A_999, A_1000;
output maj;
wire one, w0, w1, w2, w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w30, w31, w32, w33, w34, w35, w36, w37, w38, w39, w40, w41, w42, w43, w44, w45, w46, w47, w48, w49, w50, w51, w52, w53, w54, w55, w56, w57, w58, w59, w60, w61, w62, w63, w64, w65, w66, w67, w68, w69, w70, w71, w72, w73, w74, w75, w76, w77, w78, w79, w80, w81, w82, w83, w84, w85, w86, w87, w88, w89, w90, w91, w92, w93, w94, w95, w96, w97, w98, w99, w100, w101, w102, w103, w104, w105, w106, w107, w108, w109, w110, w111, w112, w113, w114, w115, w116, w117, w118, w119, w120, w121, w122, w123, w124, w125, w126, w127, w128, w129, w130, w131, w132, w133, w134, w135, w136, w137, w138, w139, w140, w141, w142, w143, w144, w145, w146, w147, w148, w149, w150, w151, w152, w153, w154, w155, w156, w157, w158, w159, w160, w161, w162, w163, w164, w165, w166, w167, w168, w169, w170, w171, w172, w173, w174, w175, w176, w177, w178, w179, w180, w181, w182, w183, w184, w185, w186, w187, w188, w189, w190, w191, w192, w193, w194, w195, w196, w197, w198, w199, w200, w201, w202, w203, w204, w205, w206, w207, w208, w209, w210, w211, w212, w213, w214, w215, w216, w217, w218, w219, w220, w221, w222, w223, w224, w225, w226, w227, w228, w229, w230, w231, w232, w233, w234, w235, w236, w237, w238, w239, w240, w241, w242, w243, w244, w245, w246, w247, w248, w249, w250, w251, w252, w253, w254, w255, w256, w257, w258, w259, w260, w261, w262, w263, w264, w265, w266, w267, w268, w269, w270, w271, w272, w273, w274, w275, w276, w277, w278, w279, w280, w281, w282, w283, w284, w285, w286, w287, w288, w289, w290, w291, w292, w293, w294, w295, w296, w297, w298, w299, w300, w301, w302, w303, w304, w305, w306, w307, w308, w309, w310, w311, w312, w313, w314, w315, w316, w317, w318, w319, w320, w321, w322, w323, w324, w325, w326, w327, w328, w329, w330, w331, w332, w333, w334, w335, w336, w337, w338, w339, w340, w341, w342, w343, w344, w345, w346, w347, w348, w349, w350, w351, w352, w353, w354, w355, w356, w357, w358, w359, w360, w361, w362, w363, w364, w365, w366, w367, w368, w369, w370, w371, w372, w373, w374, w375, w376, w377, w378, w379, w380, w381, w382, w383, w384, w385, w386, w387, w388, w389, w390, w391, w392, w393, w394, w395, w396, w397, w398, w399, w400, w401, w402, w403, w404, w405, w406, w407, w408, w409, w410, w411, w412, w413, w414, w415, w416, w417, w418, w419, w420, w421, w422, w423, w424, w425, w426, w427, w428, w429, w430, w431, w432, w433, w434, w435, w436, w437, w438, w439, w440, w441, w442, w443, w444, w445, w446, w447, w448, w449, w450, w451, w452, w453, w454, w455, w456, w457, w458, w459, w460, w461, w462, w463, w464, w465, w466, w467, w468, w469, w470, w471, w472, w473, w474, w475, w476, w477, w478, w479, w480, w481, w482, w483, w484, w485, w486, w487, w488, w489, w490, w491, w492, w493, w494, w495, w496, w497, w498, w499, w500, w501, w502, w503, w504, w505, w506, w507, w508, w509, w510, w511, w512, w513, w514, w515, w516, w517, w518, w519, w520, w521, w522, w523, w524, w525, w526, w527, w528, w529, w530, w531, w532, w533, w534, w535, w536, w537, w538, w539, w540, w541, w542, w543, w544, w545, w546, w547, w548, w549, w550, w551, w552, w553, w554, w555, w556, w557, w558, w559, w560, w561, w562, w563, w564, w565, w566, w567, w568, w569, w570, w571, w572, w573, w574, w575, w576, w577, w578, w579, w580, w581, w582, w583, w584, w585, w586, w587, w588, w589, w590, w591, w592, w593, w594, w595, w596, w597, w598, w599, w600, w601, w602, w603, w604, w605, w606, w607, w608, w609, w610, w611, w612, w613, w614, w615, w616, w617, w618, w619, w620, w621, w622, w623, w624, w625, w626, w627, w628, w629, w630, w631, w632, w633, w634, w635, w636, w637, w638, w639, w640, w641, w642, w643, w644, w645, w646, w647, w648, w649, w650, w651, w652, w653, w654, w655, w656, w657, w658, w659, w660, w661, w662, w663, w664, w665, w666, w667, w668, w669, w670, w671, w672, w673, w674, w675, w676, w677, w678, w679, w680, w681, w682, w683, w684, w685, w686, w687, w688, w689, w690, w691, w692, w693, w694, w695, w696, w697, w698, w699, w700, w701, w702, w703, w704, w705, w706, w707, w708, w709, w710, w711, w712, w713, w714, w715, w716, w717, w718, w719, w720, w721, w722, w723, w724, w725, w726, w727, w728, w729, w730, w731, w732, w733, w734, w735, w736, w737, w738, w739, w740, w741, w742, w743, w744, w745, w746, w747, w748, w749, w750, w751, w752, w753, w754, w755, w756, w757, w758, w759, w760, w761, w762, w763, w764, w765, w766, w767, w768, w769, w770, w771, w772, w773, w774, w775, w776, w777, w778, w779, w780, w781, w782, w783, w784, w785, w786, w787, w788, w789, w790, w791, w792, w793, w794, w795, w796, w797, w798, w799, w800, w801, w802, w803, w804, w805, w806, w807, w808, w809, w810, w811, w812, w813, w814, w815, w816, w817, w818, w819, w820, w821, w822, w823, w824, w825, w826, w827, w828, w829, w830, w831, w832, w833, w834, w835, w836, w837, w838, w839, w840, w841, w842, w843, w844, w845, w846, w847, w848, w849, w850, w851, w852, w853, w854, w855, w856, w857, w858, w859, w860, w861, w862, w863, w864, w865, w866, w867, w868, w869, w870, w871, w872, w873, w874, w875, w876, w877, w878, w879, w880, w881, w882, w883, w884, w885, w886, w887, w888, w889, w890, w891, w892, w893, w894, w895, w896, w897, w898, w899, w900, w901, w902, w903, w904, w905, w906, w907, w908, w909, w910, w911, w912, w913, w914, w915, w916, w917, w918, w919, w920, w921, w922, w923, w924, w925, w926, w927, w928, w929, w930, w931, w932, w933, w934, w935, w936, w937, w938, w939, w940, w941, w942, w943, w944, w945, w946, w947, w948, w949, w950, w951, w952, w953, w954, w955, w956, w957, w958, w959, w960, w961, w962, w963, w964, w965, w966, w967, w968, w969, w970, w971, w972, w973, w974, w975, w976, w977, w978, w979, w980, w981, w982, w983, w984, w985, w986, w987, w988, w989, w990, w991, w992, w993, w994, w995, w996, w997, w998, w999, w1000, w1001, w1002, w1003, w1004, w1005, w1006, w1007, w1008, w1009, w1010, w1011, w1012, w1013, w1014, w1015, w1016, w1017, w1018, w1019, w1020, w1021, w1022, w1023, w1024, w1025, w1026, w1027, w1028, w1029, w1030, w1031, w1032, w1033, w1034, w1035, w1036, w1037, w1038, w1039, w1040, w1041, w1042, w1043, w1044, w1045, w1046, w1047, w1048, w1049, w1050, w1051, w1052, w1053, w1054, w1055, w1056, w1057, w1058, w1059, w1060, w1061, w1062, w1063, w1064, w1065, w1066, w1067, w1068, w1069, w1070, w1071, w1072, w1073, w1074, w1075, w1076, w1077, w1078, w1079, w1080, w1081, w1082, w1083, w1084, w1085, w1086, w1087, w1088, w1089, w1090, w1091, w1092, w1093, w1094, w1095, w1096, w1097, w1098, w1099, w1100, w1101, w1102, w1103, w1104, w1105, w1106, w1107, w1108, w1109, w1110, w1111, w1112, w1113, w1114, w1115, w1116, w1117, w1118, w1119, w1120, w1121, w1122, w1123, w1124, w1125, w1126, w1127, w1128, w1129, w1130, w1131, w1132, w1133, w1134, w1135, w1136, w1137, w1138, w1139, w1140, w1141, w1142, w1143, w1144, w1145, w1146, w1147, w1148, w1149, w1150, w1151, w1152, w1153, w1154, w1155, w1156, w1157, w1158, w1159, w1160, w1161, w1162, w1163, w1164, w1165, w1166, w1167, w1168, w1169, w1170, w1171, w1172, w1173, w1174, w1175, w1176, w1177, w1178, w1179, w1180, w1181, w1182, w1183, w1184, w1185, w1186, w1187, w1188, w1189, w1190, w1191, w1192, w1193, w1194, w1195, w1196, w1197, w1198, w1199, w1200, w1201, w1202, w1203, w1204, w1205, w1206, w1207, w1208, w1209, w1210, w1211, w1212, w1213, w1214, w1215, w1216, w1217, w1218, w1219, w1220, w1221, w1222, w1223, w1224, w1225, w1226, w1227, w1228, w1229, w1230, w1231, w1232, w1233, w1234, w1235, w1236, w1237, w1238, w1239, w1240, w1241, w1242, w1243, w1244, w1245, w1246, w1247, w1248, w1249, w1250, w1251, w1252, w1253, w1254, w1255, w1256, w1257, w1258, w1259, w1260, w1261, w1262, w1263, w1264, w1265, w1266, w1267, w1268, w1269, w1270, w1271, w1272, w1273, w1274, w1275, w1276, w1277, w1278, w1279, w1280, w1281, w1282, w1283, w1284, w1285, w1286, w1287, w1288, w1289, w1290, w1291, w1292, w1293, w1294, w1295, w1296, w1297, w1298, w1299, w1300, w1301, w1302, w1303, w1304, w1305, w1306, w1307, w1308, w1309, w1310, w1311, w1312, w1313, w1314, w1315, w1316, w1317, w1318, w1319, w1320, w1321, w1322, w1323, w1324, w1325, w1326, w1327, w1328, w1329, w1330, w1331, w1332, w1333, w1334, w1335, w1336, w1337, w1338, w1339, w1340, w1341, w1342, w1343, w1344, w1345, w1346, w1347, w1348, w1349, w1350, w1351, w1352, w1353, w1354, w1355, w1356, w1357, w1358, w1359, w1360, w1361, w1362, w1363, w1364, w1365, w1366, w1367, w1368, w1369, w1370, w1371, w1372, w1373, w1374, w1375, w1376, w1377, w1378, w1379, w1380, w1381, w1382, w1383, w1384, w1385, w1386, w1387, w1388, w1389, w1390, w1391, w1392, w1393, w1394, w1395, w1396, w1397, w1398, w1399, w1400, w1401, w1402, w1403, w1404, w1405, w1406, w1407, w1408, w1409, w1410, w1411, w1412, w1413, w1414, w1415, w1416, w1417, w1418, w1419, w1420, w1421, w1422, w1423, w1424, w1425, w1426, w1427, w1428, w1429, w1430, w1431, w1432, w1433, w1434, w1435, w1436, w1437, w1438, w1439, w1440, w1441, w1442, w1443, w1444, w1445, w1446, w1447, w1448, w1449, w1450, w1451, w1452, w1453, w1454, w1455, w1456, w1457, w1458, w1459, w1460, w1461, w1462, w1463, w1464, w1465, w1466, w1467, w1468, w1469, w1470, w1471, w1472, w1473, w1474, w1475, w1476, w1477, w1478, w1479, w1480, w1481, w1482, w1483, w1484, w1485, w1486, w1487, w1488, w1489, w1490, w1491, w1492, w1493, w1494, w1495, w1496, w1497, w1498, w1499, w1500, w1501, w1502, w1503, w1504, w1505, w1506, w1507, w1508, w1509, w1510, w1511, w1512, w1513, w1514, w1515, w1516, w1517, w1518, w1519, w1520, w1521, w1522, w1523, w1524, w1525, w1526, w1527, w1528, w1529, w1530, w1531, w1532, w1533, w1534, w1535, w1536, w1537, w1538, w1539, w1540, w1541, w1542, w1543, w1544, w1545, w1546, w1547, w1548, w1549, w1550, w1551, w1552, w1553, w1554, w1555, w1556, w1557, w1558, w1559, w1560, w1561, w1562, w1563, w1564, w1565, w1566, w1567, w1568, w1569, w1570, w1571, w1572, w1573, w1574, w1575, w1576, w1577, w1578, w1579, w1580, w1581, w1582, w1583, w1584, w1585, w1586, w1587, w1588, w1589, w1590, w1591, w1592, w1593, w1594, w1595, w1596, w1597, w1598, w1599, w1600, w1601, w1602, w1603, w1604, w1605, w1606, w1607, w1608, w1609, w1610, w1611, w1612, w1613, w1614, w1615, w1616, w1617, w1618, w1619, w1620, w1621, w1622, w1623, w1624, w1625, w1626, w1627, w1628, w1629, w1630, w1631, w1632, w1633, w1634, w1635, w1636, w1637, w1638, w1639, w1640, w1641, w1642, w1643, w1644, w1645, w1646, w1647, w1648, w1649, w1650, w1651, w1652, w1653, w1654, w1655, w1656, w1657, w1658, w1659, w1660, w1661, w1662, w1663, w1664, w1665, w1666, w1667, w1668, w1669, w1670, w1671, w1672, w1673, w1674, w1675, w1676, w1677, w1678, w1679, w1680, w1681, w1682, w1683, w1684, w1685, w1686, w1687, w1688, w1689, w1690, w1691, w1692, w1693, w1694, w1695, w1696, w1697, w1698, w1699, w1700, w1701, w1702, w1703, w1704, w1705, w1706, w1707, w1708, w1709, w1710, w1711, w1712, w1713, w1714, w1715, w1716, w1717, w1718, w1719, w1720, w1721, w1722, w1723, w1724, w1725, w1726, w1727, w1728, w1729, w1730, w1731, w1732, w1733, w1734, w1735, w1736, w1737, w1738, w1739, w1740, w1741, w1742, w1743, w1744, w1745, w1746, w1747, w1748, w1749, w1750, w1751, w1752, w1753, w1754, w1755, w1756, w1757, w1758, w1759, w1760, w1761, w1762, w1763, w1764, w1765, w1766, w1767, w1768, w1769, w1770, w1771, w1772, w1773, w1774, w1775, w1776, w1777, w1778, w1779, w1780, w1781, w1782, w1783, w1784, w1785, w1786, w1787, w1788, w1789, w1790, w1791, w1792, w1793, w1794, w1795, w1796, w1797, w1798, w1799, w1800, w1801, w1802, w1803, w1804, w1805, w1806, w1807, w1808, w1809, w1810, w1811, w1812, w1813, w1814, w1815, w1816, w1817, w1818, w1819, w1820, w1821, w1822, w1823, w1824, w1825, w1826, w1827, w1828, w1829, w1830, w1831, w1832, w1833, w1834, w1835, w1836, w1837, w1838, w1839, w1840, w1841, w1842, w1843, w1844, w1845, w1846, w1847, w1848, w1849, w1850, w1851, w1852, w1853, w1854, w1855, w1856, w1857, w1858, w1859, w1860, w1861, w1862, w1863, w1864, w1865, w1866, w1867, w1868, w1869, w1870, w1871, w1872, w1873, w1874, w1875, w1876, w1877, w1878, w1879, w1880, w1881, w1882, w1883, w1884, w1885, w1886, w1887, w1888, w1889, w1890, w1891, w1892, w1893, w1894, w1895, w1896, w1897, w1898, w1899, w1900, w1901, w1902, w1903, w1904, w1905, w1906, w1907, w1908, w1909, w1910, w1911, w1912, w1913, w1914, w1915, w1916, w1917, w1918, w1919, w1920, w1921, w1922, w1923, w1924, w1925, w1926, w1927, w1928, w1929, w1930, w1931, w1932, w1933, w1934, w1935, w1936, w1937, w1938, w1939, w1940, w1941, w1942, w1943, w1944, w1945, w1946, w1947, w1948, w1949, w1950, w1951, w1952, w1953, w1954, w1955, w1956, w1957, w1958, w1959, w1960, w1961, w1962, w1963, w1964, w1965, w1966, w1967, w1968, w1969, w1970, w1971, w1972, w1973, w1974, w1975, w1976, w1977, w1978, w1979, w1980, w1981, w1982, w1983, w1984, w1985, w1986, w1987, w1988, w1989, w1990, w1991, w1992, w1993, w1994, w1995, w1996, w1997, w1998, w1999, w2000, w2001, w2002, w2003, w2004, w2005, w2006, w2007, w2008, w2009, w2010, w2011, w2012, w2013, w2014, w2015, w2016, w2017, w2018, w2019, w2020, w2021, w2022, w2023, w2024, w2025, w2026, w2027, w2028, w2029, w2030, w2031, w2032, w2033, w2034, w2035, w2036, w2037, w2038, w2039, w2040, w2041, w2042, w2043, w2044, w2045, w2046, w2047, w2048, w2049, w2050, w2051, w2052, w2053, w2054, w2055, w2056, w2057, w2058, w2059, w2060, w2061, w2062, w2063, w2064, w2065, w2066, w2067, w2068, w2069, w2070, w2071, w2072, w2073, w2074, w2075, w2076, w2077, w2078, w2079, w2080, w2081, w2082, w2083, w2084, w2085, w2086, w2087, w2088, w2089, w2090, w2091, w2092, w2093, w2094, w2095, w2096, w2097, w2098, w2099, w2100, w2101, w2102, w2103, w2104, w2105, w2106, w2107, w2108, w2109, w2110, w2111, w2112, w2113, w2114, w2115, w2116, w2117, w2118, w2119, w2120, w2121, w2122, w2123, w2124, w2125, w2126, w2127, w2128, w2129, w2130, w2131, w2132, w2133, w2134, w2135, w2136, w2137, w2138, w2139, w2140, w2141, w2142, w2143, w2144, w2145, w2146, w2147, w2148, w2149, w2150, w2151, w2152, w2153, w2154, w2155, w2156, w2157, w2158, w2159, w2160, w2161, w2162, w2163, w2164, w2165, w2166, w2167, w2168, w2169, w2170, w2171, w2172, w2173, w2174, w2175, w2176, w2177, w2178, w2179, w2180, w2181, w2182, w2183, w2184, w2185, w2186, w2187, w2188, w2189, w2190, w2191, w2192, w2193, w2194, w2195, w2196, w2197, w2198, w2199, w2200, w2201, w2202, w2203, w2204, w2205, w2206, w2207, w2208, w2209, w2210, w2211, w2212, w2213, w2214, w2215, w2216, w2217, w2218, w2219, w2220, w2221, w2222, w2223, w2224, w2225, w2226, w2227, w2228, w2229, w2230, w2231, w2232, w2233, w2234, w2235, w2236, w2237, w2238, w2239, w2240, w2241, w2242, w2243, w2244, w2245, w2246, w2247, w2248, w2249, w2250, w2251, w2252, w2253, w2254, w2255, w2256, w2257, w2258, w2259, w2260, w2261, w2262, w2263, w2264, w2265, w2266, w2267, w2268, w2269, w2270, w2271, w2272, w2273, w2274, w2275, w2276, w2277, w2278, w2279, w2280, w2281, w2282, w2283, w2284, w2285, w2286, w2287, w2288, w2289, w2290, w2291, w2292, w2293, w2294, w2295, w2296, w2297, w2298, w2299, w2300, w2301, w2302, w2303, w2304, w2305, w2306, w2307, w2308, w2309, w2310, w2311, w2312, w2313, w2314, w2315, w2316, w2317, w2318, w2319, w2320, w2321, w2322, w2323, w2324, w2325, w2326, w2327, w2328, w2329, w2330, w2331, w2332, w2333, w2334, w2335, w2336, w2337, w2338, w2339, w2340, w2341, w2342, w2343, w2344, w2345, w2346, w2347, w2348, w2349, w2350, w2351, w2352, w2353, w2354, w2355, w2356, w2357, w2358, w2359, w2360, w2361, w2362, w2363, w2364, w2365, w2366, w2367, w2368, w2369, w2370, w2371, w2372, w2373, w2374, w2375, w2376, w2377, w2378, w2379, w2380, w2381, w2382, w2383, w2384, w2385, w2386, w2387, w2388, w2389, w2390, w2391, w2392, w2393, w2394, w2395, w2396, w2397, w2398, w2399, w2400, w2401, w2402, w2403, w2404, w2405, w2406, w2407, w2408, w2409, w2410, w2411, w2412, w2413, w2414, w2415, w2416, w2417, w2418, w2419, w2420, w2421, w2422, w2423, w2424, w2425, w2426, w2427, w2428, w2429, w2430, w2431, w2432, w2433, w2434, w2435, w2436, w2437, w2438, w2439, w2440, w2441, w2442, w2443, w2444, w2445, w2446, w2447, w2448, w2449, w2450, w2451, w2452, w2453, w2454, w2455, w2456, w2457, w2458, w2459, w2460, w2461, w2462, w2463, w2464, w2465, w2466, w2467, w2468, w2469, w2470, w2471, w2472, w2473, w2474, w2475, w2476, w2477, w2478, w2479, w2480, w2481, w2482, w2483, w2484, w2485, w2486, w2487, w2488, w2489, w2490, w2491, w2492, w2493, w2494, w2495, w2496, w2497, w2498, w2499, w2500, w2501, w2502, w2503, w2504, w2505, w2506, w2507, w2508, w2509, w2510, w2511, w2512, w2513, w2514, w2515, w2516, w2517, w2518, w2519, w2520, w2521, w2522, w2523, w2524, w2525, w2526, w2527, w2528, w2529, w2530, w2531, w2532, w2533, w2534, w2535, w2536, w2537, w2538, w2539, w2540, w2541, w2542, w2543, w2544, w2545, w2546, w2547, w2548, w2549, w2550, w2551, w2552, w2553, w2554, w2555, w2556, w2557, w2558, w2559, w2560, w2561, w2562, w2563, w2564, w2565, w2566, w2567, w2568, w2569, w2570, w2571, w2572, w2573, w2574, w2575, w2576, w2577, w2578, w2579, w2580, w2581, w2582, w2583, w2584, w2585, w2586, w2587, w2588, w2589, w2590, w2591, w2592, w2593, w2594, w2595, w2596, w2597, w2598, w2599, w2600, w2601, w2602, w2603, w2604, w2605, w2606, w2607, w2608, w2609, w2610, w2611, w2612, w2613, w2614, w2615, w2616, w2617, w2618, w2619, w2620, w2621, w2622, w2623, w2624, w2625, w2626, w2627, w2628, w2629, w2630, w2631, w2632, w2633, w2634, w2635, w2636, w2637, w2638, w2639, w2640, w2641, w2642, w2643, w2644, w2645, w2646, w2647, w2648, w2649, w2650, w2651, w2652, w2653, w2654, w2655, w2656, w2657, w2658, w2659, w2660, w2661, w2662, w2663, w2664, w2665, w2666, w2667, w2668, w2669, w2670, w2671, w2672, w2673, w2674, w2675, w2676, w2677, w2678, w2679, w2680, w2681, w2682, w2683, w2684, w2685, w2686, w2687, w2688, w2689, w2690, w2691, w2692, w2693, w2694, w2695, w2696, w2697, w2698, w2699, w2700, w2701, w2702, w2703, w2704, w2705, w2706, w2707, w2708, w2709, w2710, w2711, w2712, w2713, w2714, w2715, w2716, w2717, w2718, w2719, w2720, w2721, w2722, w2723, w2724, w2725, w2726, w2727, w2728, w2729, w2730, w2731, w2732, w2733, w2734, w2735, w2736, w2737, w2738, w2739, w2740, w2741, w2742, w2743, w2744, w2745, w2746, w2747, w2748, w2749, w2750, w2751, w2752, w2753, w2754, w2755, w2756, w2757, w2758, w2759, w2760, w2761, w2762, w2763, w2764, w2765, w2766, w2767, w2768, w2769, w2770, w2771, w2772, w2773, w2774, w2775, w2776, w2777, w2778, w2779, w2780, w2781, w2782, w2783, w2784, w2785, w2786, w2787, w2788, w2789, w2790, w2791, w2792, w2793, w2794, w2795, w2796, w2797, w2798, w2799, w2800, w2801, w2802, w2803, w2804, w2805, w2806, w2807, w2808, w2809, w2810, w2811, w2812, w2813, w2814, w2815, w2816, w2817, w2818, w2819, w2820, w2821, w2822, w2823, w2824, w2825, w2826, w2827, w2828, w2829, w2830, w2831, w2832, w2833, w2834, w2835, w2836, w2837, w2838, w2839, w2840, w2841, w2842, w2843, w2844, w2845, w2846, w2847, w2848, w2849, w2850, w2851, w2852, w2853, w2854, w2855, w2856, w2857, w2858, w2859, w2860, w2861, w2862, w2863, w2864, w2865, w2866, w2867, w2868, w2869, w2870, w2871, w2872, w2873, w2874, w2875, w2876, w2877, w2878, w2879, w2880, w2881, w2882, w2883, w2884, w2885, w2886, w2887, w2888, w2889, w2890, w2891, w2892, w2893, w2894, w2895, w2896, w2897, w2898, w2899, w2900, w2901, w2902, w2903, w2904, w2905, w2906, w2907, w2908, w2909, w2910, w2911, w2912, w2913, w2914, w2915, w2916, w2917, w2918, w2919, w2920, w2921, w2922, w2923, w2924, w2925, w2926, w2927, w2928, w2929, w2930, w2931, w2932, w2933, w2934, w2935, w2936, w2937, w2938, w2939, w2940, w2941, w2942, w2943, w2944, w2945, w2946, w2947, w2948, w2949, w2950, w2951, w2952, w2953, w2954, w2955, w2956, w2957, w2958, w2959, w2960, w2961, w2962, w2963, w2964, w2965, w2966, w2967, w2968, w2969, w2970, w2971, w2972, w2973, w2974, w2975, w2976, w2977, w2978, w2979, w2980, w2981, w2982, w2983, w2984, w2985, w2986, w2987, w2988, w2989, w2990, w2991, w2992, w2993, w2994, w2995, w2996, w2997, w2998, w2999, w3000, w3001, w3002, w3003, w3004, w3005, w3006, w3007, w3008, w3009, w3010, w3011, w3012, w3013, w3014, w3015, w3016, w3017, w3018, w3019, w3020, w3021, w3022, w3023, w3024, w3025, w3026, w3027, w3028, w3029, w3030, w3031, w3032, w3033, w3034, w3035, w3036, w3037, w3038, w3039, w3040, w3041, w3042, w3043, w3044, w3045, w3046, w3047, w3048, w3049, w3050, w3051, w3052, w3053, w3054, w3055, w3056, w3057, w3058, w3059, w3060, w3061, w3062, w3063, w3064, w3065, w3066, w3067, w3068, w3069, w3070, w3071, w3072, w3073, w3074, w3075, w3076, w3077, w3078, w3079, w3080, w3081, w3082, w3083, w3084, w3085, w3086, w3087, w3088, w3089, w3090, w3091, w3092, w3093, w3094, w3095, w3096, w3097, w3098, w3099, w3100, w3101, w3102, w3103, w3104, w3105, w3106, w3107, w3108, w3109, w3110, w3111, w3112, w3113, w3114, w3115, w3116, w3117, w3118, w3119, w3120, w3121, w3122, w3123, w3124, w3125, w3126, w3127, w3128, w3129, w3130, w3131, w3132, w3133, w3134, w3135, w3136, w3137, w3138, w3139, w3140, w3141, w3142, w3143, w3144, w3145, w3146, w3147, w3148, w3149, w3150, w3151, w3152, w3153, w3154, w3155, w3156, w3157, w3158, w3159, w3160, w3161, w3162, w3163, w3164, w3165, w3166, w3167, w3168, w3169, w3170, w3171, w3172, w3173, w3174, w3175, w3176, w3177, w3178, w3179, w3180, w3181, w3182, w3183, w3184, w3185, w3186, w3187, w3188, w3189, w3190, w3191, w3192, w3193, w3194, w3195, w3196, w3197, w3198, w3199, w3200, w3201, w3202, w3203, w3204, w3205, w3206, w3207, w3208, w3209, w3210, w3211, w3212, w3213, w3214, w3215, w3216, w3217, w3218, w3219, w3220, w3221, w3222, w3223, w3224, w3225, w3226, w3227, w3228, w3229, w3230, w3231, w3232, w3233, w3234, w3235, w3236, w3237, w3238, w3239, w3240, w3241, w3242, w3243, w3244, w3245, w3246, w3247, w3248, w3249, w3250, w3251, w3252, w3253, w3254, w3255, w3256, w3257, w3258, w3259, w3260, w3261, w3262, w3263, w3264, w3265, w3266, w3267, w3268, w3269, w3270, w3271, w3272, w3273, w3274, w3275, w3276, w3277, w3278, w3279, w3280, w3281, w3282, w3283, w3284, w3285, w3286, w3287, w3288, w3289, w3290, w3291, w3292, w3293, w3294, w3295, w3296, w3297, w3298, w3299, w3300, w3301, w3302, w3303, w3304, w3305, w3306, w3307, w3308, w3309, w3310, w3311, w3312, w3313, w3314, w3315, w3316, w3317, w3318, w3319, w3320, w3321, w3322, w3323, w3324, w3325, w3326, w3327, w3328, w3329, w3330, w3331, w3332, w3333, w3334, w3335, w3336, w3337, w3338, w3339, w3340, w3341, w3342, w3343, w3344, w3345, w3346, w3347, w3348, w3349, w3350, w3351, w3352, w3353, w3354, w3355, w3356, w3357, w3358, w3359, w3360, w3361, w3362, w3363, w3364, w3365, w3366, w3367, w3368, w3369, w3370, w3371, w3372, w3373, w3374, w3375, w3376, w3377, w3378, w3379, w3380, w3381, w3382, w3383, w3384, w3385, w3386, w3387, w3388, w3389, w3390, w3391, w3392, w3393, w3394, w3395, w3396, w3397, w3398, w3399, w3400, w3401, w3402, w3403, w3404, w3405, w3406, w3407, w3408, w3409, w3410, w3411, w3412, w3413, w3414, w3415, w3416, w3417, w3418, w3419, w3420, w3421, w3422, w3423, w3424, w3425, w3426, w3427, w3428, w3429, w3430, w3431, w3432, w3433, w3434, w3435, w3436, w3437, w3438, w3439, w3440, w3441, w3442, w3443, w3444, w3445, w3446, w3447, w3448, w3449, w3450, w3451, w3452, w3453, w3454, w3455, w3456, w3457, w3458, w3459, w3460, w3461, w3462, w3463, w3464, w3465, w3466, w3467, w3468, w3469, w3470, w3471, w3472, w3473, w3474, w3475, w3476, w3477, w3478, w3479, w3480, w3481, w3482, w3483, w3484, w3485, w3486, w3487, w3488, w3489, w3490, w3491, w3492, w3493, w3494, w3495, w3496, w3497, w3498, w3499, w3500, w3501, w3502, w3503, w3504, w3505, w3506, w3507, w3508, w3509, w3510, w3511, w3512, w3513, w3514, w3515, w3516, w3517, w3518, w3519, w3520, w3521, w3522, w3523, w3524, w3525, w3526, w3527, w3528, w3529, w3530, w3531, w3532, w3533, w3534, w3535, w3536, w3537, w3538, w3539, w3540, w3541, w3542, w3543, w3544, w3545, w3546, w3547, w3548, w3549, w3550, w3551, w3552, w3553, w3554, w3555, w3556, w3557, w3558, w3559, w3560, w3561, w3562, w3563, w3564, w3565, w3566, w3567, w3568, w3569, w3570, w3571, w3572, w3573, w3574, w3575, w3576, w3577, w3578, w3579, w3580, w3581, w3582, w3583, w3584, w3585, w3586, w3587, w3588, w3589, w3590, w3591, w3592, w3593, w3594, w3595, w3596, w3597, w3598, w3599, w3600, w3601, w3602, w3603, w3604, w3605, w3606, w3607, w3608, w3609, w3610, w3611, w3612, w3613, w3614, w3615, w3616, w3617, w3618, w3619, w3620, w3621, w3622, w3623, w3624, w3625, w3626, w3627, w3628, w3629, w3630, w3631, w3632, w3633, w3634, w3635, w3636, w3637, w3638, w3639, w3640, w3641, w3642, w3643, w3644, w3645, w3646, w3647, w3648, w3649, w3650, w3651, w3652, w3653, w3654, w3655, w3656, w3657, w3658, w3659, w3660, w3661, w3662, w3663, w3664, w3665, w3666, w3667, w3668, w3669, w3670, w3671, w3672, w3673, w3674, w3675, w3676, w3677, w3678, w3679, w3680, w3681, w3682, w3683, w3684, w3685, w3686, w3687, w3688, w3689, w3690, w3691, w3692, w3693, w3694, w3695, w3696, w3697, w3698, w3699, w3700, w3701, w3702, w3703, w3704, w3705, w3706, w3707, w3708, w3709, w3710, w3711, w3712, w3713, w3714, w3715, w3716, w3717, w3718, w3719, w3720, w3721, w3722, w3723, w3724, w3725, w3726, w3727, w3728, w3729, w3730, w3731, w3732, w3733, w3734, w3735, w3736, w3737, w3738, w3739, w3740, w3741, w3742, w3743, w3744, w3745, w3746, w3747, w3748, w3749, w3750, w3751, w3752, w3753, w3754, w3755, w3756, w3757, w3758, w3759, w3760, w3761, w3762, w3763, w3764, w3765, w3766, w3767, w3768, w3769, w3770, w3771, w3772, w3773, w3774, w3775, w3776, w3777, w3778, w3779, w3780, w3781, w3782, w3783, w3784, w3785, w3786, w3787, w3788, w3789, w3790, w3791, w3792, w3793, w3794, w3795, w3796, w3797, w3798, w3799, w3800, w3801, w3802, w3803, w3804, w3805, w3806, w3807, w3808, w3809, w3810, w3811, w3812, w3813, w3814, w3815, w3816, w3817, w3818, w3819, w3820, w3821, w3822, w3823, w3824, w3825, w3826, w3827, w3828, w3829, w3830, w3831, w3832, w3833, w3834, w3835, w3836, w3837, w3838, w3839, w3840, w3841, w3842, w3843, w3844, w3845, w3846, w3847, w3848, w3849, w3850, w3851, w3852, w3853, w3854, w3855, w3856, w3857, w3858, w3859, w3860, w3861, w3862, w3863, w3864, w3865, w3866, w3867, w3868, w3869, w3870, w3871, w3872, w3873, w3874, w3875, w3876, w3877, w3878, w3879, w3880, w3881, w3882, w3883, w3884, w3885, w3886, w3887, w3888, w3889, w3890, w3891, w3892, w3893, w3894, w3895, w3896, w3897, w3898, w3899, w3900, w3901, w3902, w3903, w3904, w3905, w3906, w3907, w3908, w3909, w3910, w3911, w3912, w3913, w3914, w3915, w3916, w3917, w3918, w3919, w3920, w3921, w3922, w3923, w3924, w3925, w3926, w3927, w3928, w3929, w3930, w3931, w3932, w3933, w3934, w3935, w3936, w3937, w3938, w3939, w3940, w3941, w3942, w3943, w3944, w3945, w3946, w3947, w3948, w3949, w3950, w3951, w3952, w3953, w3954, w3955, w3956, w3957, w3958, w3959, w3960, w3961, w3962, w3963, w3964, w3965, w3966, w3967, w3968, w3969, w3970, w3971, w3972, w3973, w3974, w3975, w3976, w3977, w3978, w3979, w3980, w3981, w3982, w3983, w3984, w3985, w3986, w3987, w3988, w3989, w3990, w3991, w3992, w3993, w3994, w3995, w3996, w3997, w3998, w3999, w4000, w4001, w4002, w4003, w4004, w4005, w4006, w4007, w4008, w4009, w4010, w4011, w4012, w4013, w4014, w4015, w4016, w4017, w4018, w4019, w4020, w4021, w4022, w4023, w4024, w4025, w4026, w4027, w4028, w4029, w4030, w4031, w4032, w4033, w4034, w4035, w4036, w4037, w4038, w4039, w4040, w4041, w4042, w4043, w4044, w4045, w4046, w4047, w4048, w4049, w4050, w4051, w4052, w4053, w4054, w4055, w4056, w4057, w4058, w4059, w4060, w4061, w4062, w4063, w4064, w4065, w4066, w4067, w4068, w4069, w4070, w4071, w4072, w4073, w4074, w4075, w4076, w4077, w4078, w4079, w4080, w4081, w4082, w4083, w4084, w4085, w4086, w4087, w4088, w4089, w4090, w4091, w4092, w4093, w4094, w4095, w4096, w4097, w4098, w4099, w4100, w4101, w4102, w4103, w4104, w4105, w4106, w4107, w4108, w4109, w4110, w4111, w4112, w4113, w4114, w4115, w4116, w4117, w4118, w4119, w4120, w4121, w4122, w4123, w4124, w4125, w4126, w4127, w4128, w4129, w4130, w4131, w4132, w4133, w4134, w4135, w4136, w4137, w4138, w4139, w4140, w4141, w4142, w4143, w4144, w4145, w4146, w4147, w4148, w4149, w4150, w4151, w4152, w4153, w4154, w4155, w4156, w4157, w4158, w4159, w4160, w4161, w4162, w4163, w4164, w4165, w4166, w4167, w4168, w4169, w4170, w4171, w4172, w4173, w4174, w4175, w4176, w4177, w4178, w4179, w4180, w4181, w4182, w4183, w4184, w4185, w4186, w4187, w4188, w4189, w4190, w4191, w4192, w4193, w4194, w4195, w4196, w4197, w4198, w4199, w4200, w4201, w4202, w4203, w4204, w4205, w4206, w4207, w4208, w4209, w4210, w4211, w4212, w4213, w4214, w4215, w4216, w4217, w4218, w4219, w4220, w4221, w4222, w4223, w4224, w4225, w4226, w4227, w4228, w4229, w4230, w4231, w4232, w4233, w4234, w4235, w4236, w4237, w4238, w4239, w4240, w4241, w4242, w4243, w4244, w4245, w4246, w4247, w4248, w4249, w4250, w4251, w4252, w4253, w4254, w4255, w4256, w4257, w4258, w4259, w4260, w4261, w4262, w4263, w4264, w4265, w4266, w4267, w4268, w4269, w4270, w4271, w4272, w4273, w4274, w4275, w4276, w4277, w4278, w4279, w4280, w4281, w4282, w4283, w4284, w4285, w4286, w4287, w4288, w4289, w4290, w4291, w4292, w4293, w4294, w4295, w4296, w4297, w4298, w4299, w4300, w4301, w4302, w4303, w4304, w4305, w4306, w4307, w4308, w4309, w4310, w4311, w4312, w4313, w4314, w4315, w4316, w4317, w4318, w4319, w4320, w4321, w4322, w4323, w4324, w4325, w4326, w4327, w4328, w4329, w4330, w4331, w4332, w4333, w4334, w4335, w4336, w4337, w4338, w4339, w4340, w4341, w4342, w4343, w4344, w4345, w4346, w4347, w4348, w4349, w4350, w4351, w4352, w4353, w4354, w4355, w4356, w4357, w4358, w4359, w4360, w4361, w4362, w4363, w4364, w4365, w4366, w4367, w4368, w4369, w4370, w4371, w4372, w4373, w4374, w4375, w4376, w4377, w4378, w4379, w4380, w4381, w4382, w4383, w4384, w4385, w4386, w4387, w4388, w4389, w4390, w4391, w4392, w4393, w4394, w4395, w4396, w4397, w4398, w4399, w4400, w4401, w4402, w4403, w4404, w4405, w4406, w4407, w4408, w4409, w4410, w4411, w4412, w4413, w4414, w4415, w4416, w4417, w4418, w4419, w4420, w4421, w4422, w4423, w4424, w4425, w4426, w4427, w4428, w4429, w4430, w4431, w4432, w4433, w4434, w4435, w4436, w4437, w4438, w4439, w4440, w4441, w4442, w4443, w4444, w4445, w4446, w4447, w4448, w4449, w4450, w4451, w4452, w4453, w4454, w4455, w4456, w4457, w4458, w4459, w4460, w4461, w4462, w4463, w4464, w4465, w4466, w4467, w4468, w4469, w4470, w4471, w4472, w4473, w4474, w4475, w4476, w4477, w4478, w4479, w4480, w4481, w4482, w4483, w4484, w4485, w4486, w4487, w4488, w4489, w4490, w4491, w4492, w4493, w4494, w4495, w4496, w4497, w4498, w4499, w4500, w4501, w4502, w4503, w4504, w4505, w4506, w4507, w4508, w4509, w4510, w4511, w4512, w4513, w4514, w4515, w4516, w4517, w4518, w4519, w4520, w4521, w4522, w4523, w4524, w4525, w4526, w4527, w4528, w4529, w4530, w4531, w4532, w4533, w4534, w4535, w4536, w4537, w4538, w4539, w4540, w4541, w4542, w4543, w4544, w4545, w4546, w4547, w4548, w4549, w4550, w4551, w4552, w4553, w4554, w4555, w4556, w4557, w4558, w4559, w4560, w4561, w4562, w4563, w4564, w4565, w4566, w4567, w4568, w4569, w4570, w4571, w4572, w4573, w4574, w4575, w4576, w4577, w4578, w4579, w4580, w4581, w4582, w4583, w4584, w4585, w4586, w4587, w4588, w4589, w4590, w4591, w4592, w4593, w4594, w4595, w4596, w4597, w4598, w4599, w4600, w4601, w4602, w4603, w4604, w4605, w4606, w4607, w4608, w4609, w4610, w4611, w4612, w4613, w4614, w4615, w4616, w4617, w4618, w4619, w4620, w4621, w4622, w4623, w4624, w4625, w4626, w4627, w4628, w4629, w4630, w4631, w4632, w4633, w4634, w4635, w4636, w4637, w4638, w4639, w4640, w4641, w4642, w4643, w4644, w4645, w4646, w4647, w4648, w4649, w4650, w4651, w4652, w4653, w4654, w4655, w4656, w4657, w4658, w4659, w4660, w4661, w4662, w4663, w4664, w4665, w4666, w4667, w4668, w4669, w4670, w4671, w4672, w4673, w4674, w4675, w4676, w4677, w4678, w4679, w4680, w4681, w4682, w4683, w4684, w4685, w4686, w4687, w4688, w4689, w4690, w4691, w4692, w4693, w4694, w4695, w4696, w4697, w4698, w4699, w4700, w4701, w4702, w4703, w4704, w4705, w4706, w4707, w4708, w4709, w4710, w4711, w4712, w4713, w4714, w4715, w4716, w4717, w4718, w4719, w4720, w4721, w4722, w4723, w4724, w4725, w4726, w4727, w4728, w4729, w4730, w4731, w4732, w4733, w4734, w4735, w4736, w4737, w4738, w4739, w4740, w4741, w4742, w4743, w4744, w4745, w4746, w4747, w4748, w4749, w4750, w4751, w4752, w4753, w4754, w4755, w4756, w4757, w4758, w4759, w4760, w4761, w4762, w4763, w4764, w4765, w4766, w4767, w4768, w4769, w4770, w4771, w4772, w4773, w4774, w4775, w4776, w4777, w4778, w4779, w4780, w4781, w4782, w4783, w4784, w4785, w4786, w4787, w4788, w4789, w4790, w4791, w4792, w4793, w4794, w4795, w4796, w4797, w4798, w4799, w4800, w4801, w4802, w4803, w4804, w4805, w4806, w4807, w4808, w4809, w4810, w4811, w4812, w4813, w4814, w4815, w4816, w4817, w4818, w4819, w4820, w4821, w4822, w4823, w4824, w4825, w4826, w4827, w4828, w4829, w4830, w4831, w4832, w4833, w4834, w4835, w4836, w4837, w4838, w4839, w4840, w4841, w4842, w4843, w4844, w4845, w4846, w4847, w4848, w4849, w4850, w4851, w4852, w4853, w4854, w4855, w4856, w4857, w4858, w4859, w4860, w4861, w4862, w4863, w4864, w4865, w4866, w4867, w4868, w4869, w4870, w4871, w4872, w4873, w4874, w4875, w4876, w4877, w4878, w4879, w4880, w4881, w4882, w4883, w4884, w4885, w4886, w4887, w4888, w4889, w4890, w4891, w4892, w4893, w4894, w4895, w4896, w4897, w4898, w4899, w4900, w4901, w4902, w4903, w4904, w4905, w4906, w4907, w4908, w4909, w4910, w4911, w4912, w4913, w4914, w4915, w4916, w4917, w4918, w4919, w4920, w4921, w4922, w4923, w4924, w4925, w4926, w4927, w4928, w4929, w4930, w4931, w4932, w4933, w4934, w4935, w4936, w4937, w4938, w4939, w4940, w4941, w4942, w4943, w4944, w4945, w4946, w4947, w4948, w4949, w4950, w4951, w4952, w4953, w4954, w4955, w4956, w4957, w4958, w4959, w4960, w4961, w4962, w4963, w4964, w4965, w4966, w4967, w4968, w4969, w4970, w4971, w4972, w4973, w4974, w4975, w4976, w4977, w4978, w4979, w4980, w4981, w4982, w4983, w4984, w4985, w4986, w4987, w4988, w4989, w4990, w4991, w4992, w4993, w4994, w4995, w4996, w4997, w4998, w4999, w5000, w5001, w5002, w5003, w5004, w5005, w5006, w5007, w5008, w5009, w5010, w5011, w5012, w5013, w5014, w5015, w5016, w5017, w5018, w5019, w5020, w5021, w5022, w5023, w5024, w5025, w5026, w5027, w5028, w5029, w5030, w5031, w5032, w5033, w5034, w5035, w5036, w5037, w5038, w5039, w5040, w5041, w5042, w5043, w5044, w5045, w5046, w5047, w5048, w5049, w5050, w5051, w5052, w5053, w5054, w5055, w5056, w5057, w5058, w5059, w5060, w5061, w5062, w5063, w5064, w5065, w5066, w5067, w5068, w5069, w5070, w5071, w5072, w5073, w5074, w5075, w5076, w5077, w5078, w5079, w5080, w5081, w5082, w5083, w5084, w5085, w5086, w5087, w5088, w5089, w5090, w5091, w5092, w5093, w5094, w5095, w5096, w5097, w5098, w5099, w5100, w5101, w5102, w5103, w5104, w5105, w5106, w5107, w5108, w5109, w5110, w5111, w5112, w5113, w5114, w5115, w5116, w5117, w5118, w5119, w5120, w5121, w5122, w5123, w5124, w5125, w5126, w5127, w5128, w5129, w5130, w5131, w5132, w5133, w5134, w5135, w5136, w5137, w5138, w5139, w5140, w5141, w5142, w5143, w5144, w5145, w5146, w5147, w5148, w5149, w5150, w5151, w5152, w5153, w5154, w5155, w5156, w5157, w5158, w5159, w5160, w5161, w5162, w5163, w5164, w5165, w5166, w5167, w5168, w5169, w5170, w5171, w5172, w5173, w5174, w5175, w5176, w5177, w5178, w5179, w5180, w5181, w5182, w5183, w5184, w5185, w5186, w5187, w5188, w5189, w5190, w5191, w5192, w5193, w5194, w5195, w5196, w5197, w5198, w5199, w5200, w5201, w5202, w5203, w5204, w5205, w5206, w5207, w5208, w5209, w5210, w5211, w5212, w5213, w5214, w5215, w5216, w5217, w5218, w5219, w5220, w5221, w5222, w5223, w5224, w5225, w5226, w5227, w5228, w5229, w5230, w5231, w5232, w5233, w5234, w5235, w5236, w5237, w5238, w5239, w5240, w5241, w5242, w5243, w5244, w5245, w5246, w5247, w5248, w5249, w5250, w5251, w5252, w5253, w5254, w5255, w5256, w5257, w5258, w5259, w5260, w5261, w5262, w5263, w5264, w5265, w5266, w5267, w5268, w5269, w5270, w5271, w5272, w5273, w5274, w5275, w5276, w5277, w5278, w5279, w5280, w5281, w5282, w5283, w5284, w5285, w5286, w5287, w5288, w5289, w5290, w5291, w5292, w5293, w5294, w5295, w5296, w5297, w5298, w5299, w5300, w5301, w5302, w5303, w5304, w5305, w5306, w5307, w5308, w5309, w5310, w5311, w5312, w5313, w5314, w5315, w5316, w5317, w5318, w5319, w5320, w5321, w5322, w5323, w5324, w5325, w5326, w5327, w5328, w5329, w5330, w5331, w5332, w5333, w5334, w5335, w5336, w5337, w5338, w5339, w5340, w5341, w5342, w5343, w5344, w5345, w5346, w5347, w5348, w5349, w5350, w5351, w5352, w5353, w5354, w5355, w5356, w5357, w5358, w5359, w5360, w5361, w5362, w5363, w5364, w5365, w5366, w5367, w5368, w5369, w5370, w5371, w5372, w5373, w5374, w5375, w5376, w5377, w5378, w5379, w5380, w5381, w5382, w5383, w5384, w5385, w5386, w5387, w5388, w5389, w5390, w5391, w5392, w5393, w5394, w5395, w5396, w5397, w5398, w5399, w5400, w5401, w5402, w5403, w5404, w5405, w5406, w5407, w5408, w5409, w5410, w5411, w5412, w5413, w5414, w5415, w5416, w5417, w5418, w5419, w5420, w5421, w5422, w5423, w5424, w5425, w5426, w5427, w5428, w5429, w5430, w5431, w5432, w5433, w5434, w5435, w5436, w5437, w5438, w5439, w5440, w5441, w5442, w5443, w5444, w5445, w5446, w5447, w5448, w5449, w5450, w5451, w5452, w5453, w5454, w5455, w5456, w5457, w5458, w5459, w5460, w5461, w5462, w5463, w5464, w5465, w5466, w5467, w5468, w5469, w5470, w5471, w5472, w5473, w5474, w5475, w5476, w5477, w5478, w5479, w5480, w5481, w5482, w5483, w5484, w5485, w5486, w5487, w5488, w5489, w5490, w5491, w5492, w5493, w5494, w5495, w5496, w5497, w5498, w5499, w5500, w5501, w5502, w5503, w5504, w5505, w5506, w5507, w5508, w5509, w5510, w5511, w5512, w5513, w5514, w5515, w5516, w5517, w5518, w5519, w5520, w5521, w5522, w5523, w5524, w5525, w5526, w5527, w5528, w5529, w5530, w5531, w5532, w5533, w5534, w5535, w5536, w5537, w5538, w5539, w5540, w5541, w5542, w5543, w5544, w5545, w5546, w5547, w5548, w5549, w5550, w5551, w5552, w5553, w5554, w5555, w5556, w5557, w5558, w5559, w5560, w5561, w5562, w5563, w5564, w5565, w5566, w5567, w5568, w5569, w5570, w5571, w5572, w5573, w5574, w5575, w5576, w5577, w5578, w5579, w5580, w5581, w5582, w5583, w5584, w5585, w5586, w5587, w5588, w5589, w5590, w5591, w5592, w5593, w5594, w5595, w5596, w5597, w5598, w5599, w5600, w5601, w5602, w5603, w5604, w5605, w5606, w5607, w5608, w5609, w5610, w5611, w5612, w5613, w5614, w5615, w5616, w5617, w5618, w5619, w5620, w5621, w5622, w5623, w5624, w5625, w5626, w5627, w5628, w5629, w5630, w5631, w5632, w5633, w5634, w5635, w5636, w5637, w5638, w5639, w5640, w5641, w5642, w5643, w5644, w5645, w5646, w5647, w5648, w5649, w5650, w5651, w5652, w5653, w5654, w5655, w5656, w5657, w5658, w5659, w5660, w5661, w5662, w5663, w5664, w5665, w5666, w5667, w5668, w5669, w5670, w5671, w5672, w5673, w5674, w5675, w5676, w5677, w5678, w5679, w5680, w5681, w5682, w5683, w5684, w5685, w5686, w5687, w5688, w5689, w5690, w5691, w5692, w5693, w5694, w5695, w5696, w5697, w5698, w5699, w5700, w5701, w5702, w5703, w5704, w5705, w5706, w5707, w5708, w5709, w5710, w5711, w5712, w5713, w5714, w5715, w5716, w5717, w5718, w5719, w5720, w5721, w5722, w5723, w5724, w5725, w5726, w5727, w5728, w5729, w5730, w5731, w5732, w5733, w5734, w5735, w5736, w5737, w5738, w5739, w5740, w5741, w5742, w5743, w5744, w5745, w5746, w5747, w5748, w5749, w5750, w5751, w5752, w5753, w5754, w5755, w5756, w5757, w5758, w5759, w5760, w5761, w5762, w5763, w5764, w5765, w5766, w5767, w5768, w5769, w5770, w5771, w5772, w5773, w5774, w5775, w5776, w5777, w5778, w5779, w5780, w5781, w5782, w5783, w5784, w5785, w5786, w5787, w5788, w5789, w5790, w5791, w5792, w5793, w5794, w5795, w5796, w5797, w5798, w5799, w5800, w5801, w5802, w5803, w5804, w5805, w5806, w5807, w5808, w5809, w5810, w5811, w5812, w5813, w5814, w5815, w5816, w5817, w5818, w5819, w5820, w5821, w5822, w5823, w5824, w5825, w5826, w5827, w5828, w5829, w5830, w5831, w5832, w5833, w5834, w5835, w5836, w5837, w5838, w5839, w5840, w5841, w5842, w5843, w5844, w5845, w5846, w5847, w5848, w5849, w5850, w5851, w5852, w5853, w5854, w5855, w5856, w5857, w5858, w5859, w5860, w5861, w5862, w5863, w5864, w5865, w5866, w5867, w5868, w5869, w5870, w5871, w5872, w5873, w5874, w5875, w5876, w5877, w5878, w5879, w5880, w5881, w5882, w5883, w5884, w5885, w5886, w5887, w5888, w5889, w5890, w5891, w5892, w5893, w5894, w5895, w5896, w5897, w5898, w5899, w5900, w5901, w5902, w5903, w5904, w5905, w5906, w5907, w5908, w5909, w5910, w5911, w5912, w5913, w5914, w5915, w5916, w5917, w5918, w5919, w5920, w5921, w5922, w5923, w5924, w5925, w5926, w5927, w5928, w5929, w5930, w5931, w5932, w5933, w5934, w5935, w5936, w5937, w5938, w5939, w5940, w5941, w5942, w5943, w5944, w5945, w5946, w5947, w5948, w5949, w5950, w5951, w5952, w5953, w5954, w5955, w5956, w5957, w5958, w5959, w5960, w5961, w5962, w5963, w5964, w5965, w5966, w5967, w5968, w5969, w5970, w5971, w5972, w5973, w5974, w5975, w5976, w5977, w5978, w5979, w5980, w5981, w5982, w5983, w5984, w5985, w5986, w5987, w5988, w5989, w5990, w5991, w5992, w5993, w5994, w5995, w5996, w5997, w5998, w5999, w6000, w6001, w6002, w6003, w6004, w6005, w6006, w6007, w6008, w6009, w6010, w6011, w6012, w6013, w6014, w6015, w6016, w6017, w6018, w6019, w6020, w6021, w6022, w6023, w6024, w6025, w6026, w6027, w6028, w6029, w6030, w6031, w6032, w6033, w6034, w6035, w6036, w6037, w6038, w6039, w6040, w6041, w6042, w6043, w6044, w6045, w6046, w6047, w6048, w6049, w6050, w6051, w6052, w6053, w6054, w6055, w6056, w6057, w6058, w6059, w6060, w6061, w6062, w6063, w6064, w6065, w6066, w6067, w6068, w6069, w6070, w6071, w6072, w6073, w6074, w6075, w6076, w6077, w6078, w6079, w6080, w6081, w6082, w6083, w6084, w6085, w6086, w6087, w6088, w6089, w6090, w6091, w6092, w6093, w6094, w6095, w6096, w6097, w6098, w6099, w6100, w6101, w6102, w6103, w6104, w6105, w6106, w6107, w6108, w6109, w6110, w6111, w6112, w6113, w6114, w6115, w6116, w6117, w6118, w6119, w6120, w6121, w6122, w6123, w6124, w6125, w6126, w6127, w6128, w6129, w6130, w6131, w6132, w6133, w6134, w6135, w6136, w6137, w6138, w6139, w6140, w6141, w6142, w6143, w6144, w6145, w6146, w6147, w6148, w6149, w6150, w6151, w6152, w6153, w6154, w6155, w6156, w6157, w6158, w6159, w6160, w6161, w6162, w6163, w6164, w6165, w6166, w6167, w6168, w6169, w6170, w6171, w6172, w6173, w6174, w6175, w6176, w6177, w6178, w6179, w6180, w6181, w6182, w6183, w6184, w6185, w6186, w6187, w6188, w6189, w6190, w6191, w6192, w6193, w6194, w6195, w6196, w6197, w6198, w6199, w6200, w6201, w6202, w6203, w6204, w6205, w6206, w6207, w6208, w6209, w6210, w6211, w6212, w6213, w6214, w6215, w6216, w6217, w6218, w6219, w6220, w6221, w6222, w6223, w6224, w6225, w6226, w6227, w6228, w6229, w6230, w6231, w6232, w6233, w6234, w6235, w6236, w6237, w6238, w6239, w6240, w6241, w6242, w6243, w6244, w6245, w6246, w6247, w6248, w6249, w6250, w6251, w6252, w6253, w6254, w6255, w6256, w6257, w6258, w6259, w6260, w6261, w6262, w6263, w6264, w6265, w6266, w6267, w6268, w6269, w6270, w6271, w6272, w6273, w6274, w6275, w6276, w6277, w6278, w6279, w6280, w6281, w6282, w6283, w6284, w6285, w6286, w6287, w6288, w6289, w6290, w6291, w6292, w6293, w6294, w6295, w6296, w6297, w6298, w6299, w6300, w6301, w6302, w6303, w6304, w6305, w6306, w6307, w6308, w6309, w6310, w6311, w6312, w6313, w6314, w6315, w6316, w6317, w6318, w6319, w6320, w6321, w6322, w6323, w6324, w6325, w6326, w6327, w6328, w6329, w6330, w6331, w6332, w6333, w6334, w6335, w6336, w6337, w6338, w6339, w6340, w6341, w6342, w6343, w6344, w6345, w6346, w6347, w6348, w6349, w6350, w6351, w6352, w6353, w6354, w6355, w6356, w6357, w6358, w6359, w6360, w6361, w6362, w6363, w6364, w6365, w6366, w6367, w6368, w6369, w6370, w6371, w6372, w6373, w6374, w6375, w6376, w6377, w6378, w6379, w6380, w6381, w6382, w6383, w6384, w6385, w6386, w6387, w6388, w6389, w6390, w6391, w6392, w6393, w6394, w6395, w6396, w6397, w6398, w6399, w6400, w6401, w6402, w6403, w6404, w6405, w6406, w6407, w6408, w6409, w6410, w6411, w6412, w6413, w6414, w6415, w6416, w6417, w6418, w6419, w6420, w6421, w6422, w6423, w6424, w6425, w6426, w6427, w6428, w6429, w6430, w6431, w6432, w6433, w6434, w6435, w6436, w6437, w6438, w6439, w6440, w6441, w6442, w6443, w6444, w6445, w6446, w6447, w6448, w6449, w6450, w6451, w6452, w6453, w6454, w6455, w6456, w6457, w6458, w6459, w6460, w6461, w6462, w6463, w6464, w6465, w6466, w6467, w6468, w6469, w6470, w6471, w6472, w6473, w6474, w6475, w6476, w6477, w6478, w6479, w6480, w6481, w6482, w6483, w6484, w6485, w6486, w6487, w6488, w6489, w6490, w6491, w6492, w6493, w6494, w6495, w6496, w6497, w6498, w6499, w6500, w6501, w6502, w6503, w6504, w6505, w6506, w6507, w6508, w6509, w6510, w6511, w6512, w6513, w6514, w6515, w6516, w6517, w6518, w6519, w6520, w6521, w6522, w6523, w6524, w6525, w6526, w6527, w6528, w6529, w6530, w6531, w6532, w6533, w6534, w6535, w6536, w6537, w6538, w6539, w6540, w6541, w6542, w6543, w6544, w6545, w6546, w6547, w6548, w6549, w6550, w6551, w6552, w6553, w6554, w6555, w6556, w6557, w6558, w6559, w6560, w6561, w6562, w6563, w6564, w6565, w6566, w6567, w6568, w6569, w6570, w6571, w6572, w6573, w6574, w6575, w6576, w6577, w6578, w6579, w6580, w6581, w6582, w6583, w6584, w6585, w6586, w6587, w6588, w6589, w6590, w6591, w6592, w6593, w6594, w6595, w6596, w6597, w6598, w6599, w6600, w6601, w6602, w6603, w6604, w6605, w6606, w6607, w6608, w6609, w6610, w6611, w6612, w6613, w6614, w6615, w6616, w6617, w6618, w6619, w6620, w6621, w6622, w6623, w6624, w6625, w6626, w6627, w6628, w6629, w6630, w6631, w6632, w6633, w6634, w6635, w6636, w6637, w6638, w6639, w6640, w6641, w6642, w6643, w6644, w6645, w6646, w6647, w6648, w6649, w6650, w6651, w6652, w6653, w6654, w6655, w6656, w6657, w6658, w6659, w6660, w6661, w6662, w6663, w6664, w6665, w6666, w6667, w6668, w6669, w6670, w6671, w6672, w6673, w6674, w6675, w6676, w6677, w6678, w6679, w6680, w6681, w6682, w6683, w6684, w6685, w6686, w6687, w6688, w6689, w6690, w6691, w6692, w6693, w6694, w6695, w6696, w6697, w6698, w6699, w6700, w6701, w6702, w6703, w6704, w6705, w6706, w6707, w6708, w6709, w6710, w6711, w6712, w6713, w6714, w6715, w6716, w6717, w6718, w6719, w6720, w6721, w6722, w6723, w6724, w6725, w6726, w6727, w6728, w6729, w6730, w6731, w6732, w6733, w6734, w6735, w6736, w6737, w6738, w6739, w6740, w6741, w6742, w6743, w6744, w6745, w6746, w6747, w6748, w6749, w6750, w6751, w6752, w6753, w6754, w6755, w6756, w6757, w6758, w6759, w6760, w6761, w6762, w6763, w6764, w6765, w6766, w6767, w6768, w6769, w6770, w6771, w6772, w6773, w6774, w6775, w6776, w6777, w6778, w6779, w6780, w6781, w6782, w6783, w6784, w6785, w6786, w6787, w6788, w6789, w6790, w6791, w6792, w6793, w6794, w6795, w6796, w6797, w6798, w6799, w6800, w6801, w6802, w6803, w6804, w6805, w6806, w6807, w6808, w6809, w6810, w6811, w6812, w6813, w6814, w6815, w6816, w6817, w6818, w6819, w6820, w6821, w6822, w6823, w6824, w6825, w6826, w6827, w6828, w6829, w6830, w6831, w6832, w6833, w6834, w6835, w6836, w6837, w6838, w6839, w6840, w6841, w6842, w6843, w6844, w6845, w6846, w6847, w6848, w6849, w6850, w6851, w6852, w6853, w6854, w6855, w6856, w6857, w6858, w6859, w6860, w6861, w6862, w6863, w6864, w6865, w6866, w6867, w6868, w6869, w6870, w6871, w6872, w6873, w6874, w6875, w6876, w6877, w6878, w6879, w6880, w6881, w6882, w6883, w6884, w6885, w6886, w6887, w6888, w6889, w6890, w6891, w6892, w6893, w6894, w6895, w6896, w6897, w6898, w6899, w6900, w6901, w6902, w6903, w6904, w6905, w6906, w6907, w6908, w6909, w6910, w6911, w6912, w6913, w6914, w6915, w6916, w6917, w6918, w6919, w6920, w6921, w6922, w6923, w6924, w6925, w6926, w6927, w6928, w6929, w6930, w6931, w6932, w6933, w6934, w6935, w6936, w6937, w6938, w6939, w6940, w6941, w6942, w6943, w6944, w6945, w6946, w6947, w6948, w6949, w6950, w6951, w6952, w6953, w6954, w6955, w6956, w6957, w6958, w6959, w6960, w6961, w6962, w6963, w6964, w6965, w6966, w6967, w6968, w6969, w6970, w6971, w6972, w6973, w6974, w6975, w6976, w6977, w6978, w6979, w6980, w6981, w6982, w6983, w6984, w6985, w6986, w6987, w6988, w6989, w6990, w6991, w6992, w6993, w6994, w6995, w6996, w6997, w6998, w6999, w7000, w7001, w7002, w7003, w7004, w7005, w7006, w7007, w7008, w7009, w7010, w7011, w7012, w7013, w7014, w7015, w7016, w7017, w7018, w7019, w7020, w7021, w7022, w7023, w7024, w7025, w7026, w7027, w7028, w7029, w7030, w7031, w7032, w7033, w7034, w7035, w7036, w7037, w7038, w7039, w7040, w7041, w7042, w7043, w7044, w7045, w7046, w7047, w7048, w7049, w7050, w7051, w7052, w7053, w7054, w7055, w7056, w7057, w7058, w7059, w7060, w7061, w7062, w7063, w7064, w7065, w7066, w7067, w7068, w7069, w7070, w7071, w7072, w7073, w7074, w7075, w7076, w7077, w7078, w7079, w7080, w7081, w7082, w7083, w7084, w7085, w7086, w7087, w7088, w7089, w7090, w7091, w7092, w7093, w7094, w7095, w7096, w7097, w7098, w7099, w7100, w7101, w7102, w7103, w7104, w7105, w7106, w7107, w7108, w7109, w7110, w7111, w7112, w7113, w7114, w7115, w7116, w7117, w7118, w7119, w7120, w7121, w7122, w7123, w7124, w7125, w7126, w7127, w7128, w7129, w7130, w7131, w7132, w7133, w7134, w7135, w7136, w7137, w7138, w7139, w7140, w7141, w7142, w7143, w7144, w7145, w7146, w7147, w7148, w7149, w7150, w7151, w7152, w7153, w7154, w7155, w7156, w7157, w7158, w7159, w7160, w7161, w7162, w7163, w7164, w7165, w7166, w7167, w7168, w7169, w7170, w7171, w7172, w7173, w7174, w7175, w7176, w7177, w7178, w7179, w7180, w7181, w7182, w7183, w7184, w7185, w7186, w7187, w7188, w7189, w7190, w7191, w7192, w7193, w7194, w7195, w7196, w7197, w7198, w7199, w7200, w7201, w7202, w7203, w7204, w7205, w7206, w7207, w7208, w7209, w7210, w7211, w7212, w7213, w7214, w7215, w7216, w7217, w7218, w7219, w7220, w7221, w7222, w7223, w7224, w7225, w7226, w7227, w7228, w7229, w7230, w7231, w7232, w7233, w7234, w7235, w7236, w7237, w7238, w7239, w7240, w7241, w7242, w7243, w7244, w7245, w7246, w7247, w7248, w7249, w7250, w7251, w7252, w7253, w7254, w7255, w7256, w7257, w7258, w7259, w7260, w7261, w7262, w7263, w7264, w7265, w7266, w7267, w7268, w7269, w7270, w7271, w7272, w7273, w7274, w7275, w7276, w7277, w7278, w7279, w7280, w7281, w7282, w7283, w7284, w7285, w7286, w7287, w7288, w7289, w7290, w7291, w7292, w7293, w7294, w7295, w7296, w7297, w7298, w7299, w7300, w7301, w7302, w7303, w7304, w7305, w7306, w7307, w7308, w7309, w7310, w7311, w7312, w7313, w7314, w7315, w7316, w7317, w7318, w7319, w7320, w7321, w7322, w7323, w7324, w7325, w7326, w7327, w7328, w7329, w7330, w7331, w7332, w7333, w7334, w7335, w7336, w7337, w7338, w7339, w7340, w7341, w7342, w7343, w7344, w7345, w7346, w7347, w7348, w7349, w7350, w7351, w7352, w7353, w7354, w7355, w7356, w7357, w7358, w7359, w7360, w7361, w7362, w7363, w7364, w7365, w7366, w7367, w7368, w7369, w7370, w7371, w7372, w7373, w7374, w7375, w7376, w7377, w7378, w7379, w7380, w7381, w7382, w7383, w7384, w7385, w7386, w7387, w7388, w7389, w7390, w7391, w7392, w7393, w7394, w7395, w7396, w7397, w7398, w7399, w7400, w7401, w7402, w7403, w7404, w7405, w7406, w7407, w7408, w7409, w7410, w7411, w7412, w7413, w7414, w7415, w7416, w7417, w7418, w7419, w7420, w7421, w7422, w7423, w7424, w7425, w7426, w7427, w7428, w7429, w7430, w7431, w7432, w7433, w7434, w7435, w7436, w7437, w7438, w7439, w7440, w7441, w7442, w7443, w7444, w7445, w7446, w7447, w7448, w7449, w7450, w7451, w7452, w7453, w7454, w7455, w7456, w7457, w7458, w7459, w7460, w7461, w7462, w7463, w7464, w7465, w7466, w7467, w7468, w7469, w7470, w7471, w7472, w7473, w7474, w7475, w7476, w7477, w7478, w7479, w7480, w7481, w7482, w7483, w7484, w7485, w7486, w7487, w7488, w7489, w7490, w7491, w7492, w7493, w7494, w7495, w7496, w7497, w7498, w7499, w7500, w7501, w7502, w7503, w7504, w7505, w7506, w7507, w7508, w7509, w7510, w7511, w7512, w7513, w7514, w7515, w7516, w7517, w7518, w7519, w7520, w7521, w7522, w7523, w7524, w7525, w7526, w7527, w7528, w7529, w7530, w7531, w7532, w7533, w7534, w7535, w7536, w7537, w7538, w7539, w7540, w7541, w7542, w7543, w7544, w7545, w7546, w7547, w7548, w7549, w7550, w7551, w7552, w7553, w7554, w7555, w7556, w7557, w7558, w7559, w7560, w7561, w7562, w7563, w7564, w7565, w7566, w7567, w7568, w7569, w7570, w7571, w7572, w7573, w7574, w7575, w7576, w7577, w7578, w7579, w7580, w7581, w7582, w7583, w7584, w7585, w7586, w7587, w7588, w7589, w7590, w7591, w7592, w7593, w7594, w7595, w7596, w7597, w7598, w7599, w7600, w7601, w7602, w7603, w7604, w7605, w7606, w7607, w7608, w7609, w7610, w7611, w7612, w7613, w7614, w7615, w7616, w7617, w7618, w7619, w7620, w7621, w7622, w7623, w7624, w7625, w7626, w7627, w7628, w7629, w7630, w7631, w7632, w7633, w7634, w7635, w7636, w7637, w7638, w7639, w7640, w7641, w7642, w7643, w7644, w7645, w7646, w7647, w7648, w7649, w7650, w7651, w7652, w7653, w7654, w7655, w7656, w7657, w7658, w7659, w7660, w7661, w7662, w7663, w7664, w7665, w7666, w7667, w7668, w7669, w7670, w7671, w7672, w7673, w7674, w7675, w7676, w7677, w7678, w7679, w7680, w7681, w7682, w7683, w7684, w7685, w7686, w7687, w7688, w7689, w7690, w7691, w7692, w7693, w7694, w7695, w7696, w7697, w7698, w7699, w7700, w7701, w7702, w7703, w7704, w7705, w7706, w7707, w7708, w7709, w7710, w7711, w7712, w7713, w7714, w7715, w7716, w7717, w7718, w7719, w7720, w7721, w7722, w7723, w7724, w7725, w7726, w7727, w7728, w7729, w7730, w7731, w7732, w7733, w7734, w7735, w7736, w7737, w7738, w7739, w7740, w7741, w7742, w7743, w7744, w7745, w7746, w7747, w7748, w7749, w7750, w7751, w7752, w7753, w7754, w7755, w7756, w7757, w7758, w7759, w7760, w7761, w7762, w7763, w7764, w7765, w7766, w7767, w7768, w7769, w7770, w7771, w7772, w7773, w7774, w7775, w7776, w7777, w7778, w7779, w7780, w7781, w7782, w7783, w7784, w7785, w7786, w7787, w7788, w7789, w7790, w7791, w7792, w7793, w7794, w7795, w7796, w7797, w7798, w7799, w7800, w7801, w7802, w7803, w7804, w7805, w7806, w7807, w7808, w7809, w7810, w7811, w7812, w7813, w7814, w7815, w7816, w7817, w7818, w7819, w7820, w7821, w7822, w7823, w7824, w7825, w7826, w7827, w7828, w7829, w7830, w7831, w7832, w7833, w7834, w7835, w7836, w7837, w7838, w7839, w7840, w7841, w7842, w7843, w7844, w7845, w7846, w7847, w7848, w7849, w7850, w7851, w7852, w7853, w7854, w7855, w7856, w7857, w7858, w7859, w7860, w7861, w7862, w7863, w7864, w7865, w7866, w7867, w7868, w7869, w7870, w7871, w7872, w7873, w7874, w7875, w7876, w7877, w7878, w7879, w7880, w7881, w7882, w7883, w7884, w7885, w7886, w7887, w7888, w7889, w7890, w7891, w7892, w7893, w7894, w7895, w7896, w7897, w7898, w7899, w7900, w7901, w7902, w7903, w7904, w7905, w7906, w7907, w7908, w7909, w7910, w7911, w7912, w7913, w7914, w7915, w7916, w7917, w7918, w7919, w7920, w7921, w7922, w7923, w7924, w7925, w7926, w7927, w7928, w7929, w7930, w7931, w7932, w7933, w7934, w7935, w7936, w7937, w7938, w7939, w7940, w7941, w7942, w7943, w7944, w7945, w7946, w7947, w7948, w7949, w7950, w7951, w7952, w7953, w7954, w7955, w7956, w7957, w7958, w7959, w7960, w7961, w7962, w7963, w7964, w7965, w7966, w7967, w7968, w7969, w7970, w7971, w7972, w7973, w7974, w7975, w7976, w7977, w7978, w7979, w7980, w7981, w7982, w7983, w7984, w7985, w7986, w7987, w7988, w7989, w7990, w7991, w7992, w7993, w7994, w7995, w7996, w7997, w7998, w7999, w8000, w8001, w8002, w8003, w8004, w8005, w8006, w8007, w8008, w8009, w8010, w8011, w8012, w8013, w8014, w8015, w8016, w8017, w8018, w8019, w8020, w8021, w8022, w8023, w8024, w8025, w8026, w8027, w8028, w8029, w8030, w8031, w8032, w8033, w8034, w8035, w8036, w8037, w8038, w8039, w8040, w8041, w8042, w8043, w8044, w8045, w8046, w8047, w8048, w8049, w8050, w8051, w8052, w8053, w8054, w8055, w8056, w8057, w8058, w8059, w8060, w8061, w8062, w8063, w8064, w8065, w8066, w8067, w8068, w8069, w8070, w8071, w8072, w8073, w8074, w8075, w8076, w8077, w8078, w8079, w8080, w8081, w8082, w8083, w8084, w8085, w8086, w8087, w8088, w8089, w8090, w8091, w8092, w8093, w8094, w8095, w8096, w8097, w8098, w8099, w8100, w8101, w8102, w8103, w8104, w8105, w8106, w8107, w8108, w8109, w8110, w8111, w8112, w8113, w8114, w8115, w8116, w8117, w8118, w8119, w8120, w8121, w8122, w8123, w8124, w8125, w8126, w8127, w8128, w8129, w8130, w8131, w8132, w8133, w8134, w8135, w8136, w8137, w8138, w8139, w8140, w8141, w8142, w8143, w8144, w8145, w8146, w8147, w8148, w8149, w8150, w8151, w8152, w8153, w8154, w8155, w8156, w8157, w8158, w8159, w8160, w8161, w8162, w8163, w8164, w8165, w8166, w8167, w8168, w8169, w8170, w8171, w8172, w8173, w8174, w8175, w8176, w8177, w8178, w8179, w8180, w8181, w8182, w8183, w8184, w8185, w8186, w8187, w8188, w8189, w8190, w8191, w8192, w8193, w8194, w8195, w8196, w8197, w8198, w8199, w8200, w8201, w8202, w8203, w8204, w8205, w8206, w8207, w8208, w8209, w8210, w8211, w8212, w8213, w8214, w8215, w8216, w8217, w8218, w8219, w8220, w8221, w8222, w8223, w8224, w8225, w8226, w8227, w8228, w8229, w8230, w8231, w8232, w8233, w8234, w8235, w8236, w8237, w8238, w8239, w8240, w8241, w8242, w8243, w8244, w8245, w8246, w8247, w8248, w8249, w8250, w8251, w8252, w8253, w8254, w8255, w8256, w8257, w8258, w8259, w8260, w8261, w8262, w8263, w8264, w8265, w8266, w8267, w8268, w8269, w8270, w8271, w8272, w8273, w8274, w8275, w8276, w8277, w8278, w8279, w8280, w8281, w8282, w8283, w8284, w8285, w8286, w8287, w8288, w8289, w8290, w8291, w8292, w8293, w8294, w8295, w8296, w8297, w8298, w8299, w8300, w8301, w8302, w8303, w8304, w8305, w8306, w8307, w8308, w8309, w8310, w8311, w8312, w8313, w8314, w8315, w8316, w8317, w8318, w8319, w8320, w8321, w8322, w8323, w8324, w8325, w8326, w8327, w8328, w8329, w8330, w8331, w8332, w8333, w8334, w8335, w8336, w8337, w8338, w8339, w8340, w8341, w8342, w8343, w8344, w8345, w8346, w8347, w8348, w8349, w8350, w8351, w8352, w8353, w8354, w8355, w8356, w8357, w8358, w8359, w8360, w8361, w8362, w8363, w8364, w8365, w8366, w8367, w8368, w8369, w8370, w8371, w8372, w8373, w8374, w8375, w8376, w8377, w8378, w8379, w8380, w8381, w8382, w8383, w8384, w8385, w8386, w8387, w8388, w8389, w8390, w8391, w8392, w8393, w8394, w8395, w8396, w8397, w8398, w8399, w8400, w8401, w8402, w8403, w8404, w8405, w8406, w8407, w8408, w8409, w8410, w8411, w8412, w8413, w8414, w8415, w8416, w8417, w8418, w8419, w8420, w8421, w8422, w8423, w8424, w8425, w8426, w8427, w8428, w8429, w8430, w8431, w8432, w8433, w8434, w8435, w8436, w8437, w8438, w8439, w8440, w8441, w8442, w8443, w8444, w8445, w8446, w8447, w8448, w8449, w8450, w8451, w8452, w8453, w8454, w8455, w8456, w8457, w8458, w8459, w8460, w8461, w8462, w8463, w8464, w8465, w8466, w8467, w8468, w8469, w8470, w8471, w8472, w8473, w8474, w8475, w8476, w8477, w8478, w8479, w8480, w8481, w8482, w8483, w8484, w8485, w8486, w8487, w8488, w8489, w8490, w8491, w8492, w8493, w8494, w8495, w8496, w8497, w8498, w8499, w8500, w8501, w8502, w8503, w8504, w8505, w8506, w8507, w8508, w8509, w8510, w8511, w8512, w8513, w8514, w8515, w8516, w8517, w8518, w8519, w8520, w8521, w8522, w8523, w8524, w8525, w8526, w8527, w8528, w8529, w8530, w8531, w8532, w8533, w8534, w8535, w8536, w8537, w8538, w8539, w8540, w8541, w8542, w8543, w8544, w8545, w8546, w8547, w8548, w8549, w8550, w8551, w8552, w8553, w8554, w8555, w8556, w8557, w8558, w8559, w8560, w8561, w8562, w8563, w8564, w8565, w8566, w8567, w8568, w8569, w8570, w8571, w8572, w8573, w8574, w8575, w8576, w8577, w8578, w8579, w8580, w8581, w8582, w8583, w8584, w8585, w8586, w8587, w8588, w8589, w8590, w8591, w8592, w8593, w8594, w8595, w8596, w8597, w8598, w8599, w8600, w8601, w8602, w8603, w8604, w8605, w8606, w8607, w8608, w8609, w8610, w8611, w8612, w8613, w8614, w8615, w8616, w8617, w8618, w8619, w8620, w8621, w8622, w8623, w8624, w8625, w8626, w8627, w8628, w8629, w8630, w8631, w8632, w8633, w8634, w8635, w8636, w8637, w8638, w8639, w8640, w8641, w8642, w8643, w8644, w8645, w8646, w8647, w8648, w8649, w8650, w8651, w8652, w8653, w8654, w8655, w8656, w8657, w8658, w8659, w8660, w8661, w8662, w8663, w8664, w8665, w8666, w8667, w8668, w8669, w8670, w8671, w8672, w8673, w8674, w8675, w8676, w8677, w8678, w8679, w8680, w8681, w8682, w8683, w8684, w8685, w8686, w8687, w8688, w8689, w8690, w8691, w8692, w8693, w8694, w8695, w8696, w8697, w8698, w8699, w8700, w8701, w8702, w8703, w8704, w8705, w8706, w8707, w8708, w8709, w8710, w8711, w8712, w8713, w8714, w8715, w8716, w8717, w8718, w8719, w8720, w8721, w8722, w8723, w8724, w8725, w8726, w8727, w8728, w8729, w8730, w8731, w8732, w8733, w8734, w8735, w8736, w8737, w8738, w8739, w8740, w8741, w8742, w8743, w8744, w8745, w8746, w8747, w8748, w8749, w8750, w8751, w8752, w8753, w8754, w8755, w8756, w8757, w8758, w8759, w8760, w8761, w8762, w8763, w8764, w8765, w8766, w8767, w8768, w8769, w8770, w8771, w8772, w8773, w8774, w8775, w8776, w8777, w8778, w8779, w8780, w8781, w8782, w8783, w8784, w8785, w8786, w8787, w8788, w8789, w8790, w8791, w8792, w8793, w8794, w8795, w8796, w8797, w8798, w8799, w8800, w8801, w8802, w8803, w8804, w8805, w8806, w8807, w8808, w8809, w8810, w8811, w8812, w8813, w8814, w8815, w8816, w8817, w8818, w8819, w8820, w8821, w8822, w8823, w8824, w8825, w8826, w8827, w8828, w8829, w8830, w8831, w8832, w8833, w8834, w8835, w8836, w8837, w8838, w8839, w8840, w8841, w8842, w8843, w8844, w8845, w8846, w8847, w8848, w8849, w8850, w8851, w8852, w8853, w8854, w8855, w8856, w8857, w8858, w8859, w8860, w8861, w8862, w8863, w8864, w8865, w8866, w8867, w8868, w8869, w8870, w8871, w8872, w8873, w8874, w8875, w8876, w8877, w8878, w8879, w8880, w8881, w8882, w8883, w8884, w8885, w8886, w8887, w8888, w8889, w8890, w8891, w8892, w8893, w8894, w8895, w8896, w8897, w8898, w8899, w8900, w8901, w8902, w8903, w8904, w8905, w8906, w8907, w8908, w8909, w8910, w8911, w8912, w8913, w8914, w8915, w8916, w8917, w8918, w8919, w8920, w8921, w8922, w8923, w8924, w8925, w8926, w8927, w8928, w8929, w8930, w8931, w8932, w8933, w8934, w8935, w8936, w8937, w8938, w8939, w8940, w8941, w8942, w8943, w8944, w8945, w8946, w8947, w8948, w8949, w8950, w8951, w8952, w8953, w8954, w8955, w8956, w8957, w8958, w8959, w8960, w8961, w8962, w8963, w8964, w8965, w8966, w8967, w8968, w8969, w8970, w8971, w8972, w8973, w8974, w8975, w8976, w8977, w8978, w8979, w8980, w8981, w8982, w8983, w8984, w8985, w8986, w8987, w8988, w8989, w8990, w8991, w8992, w8993, w8994, w8995, w8996, w8997, w8998, w8999, w9000, w9001, w9002, w9003, w9004, w9005, w9006, w9007, w9008, w9009, w9010, w9011, w9012, w9013, w9014, w9015, w9016, w9017, w9018, w9019, w9020, w9021, w9022, w9023, w9024, w9025, w9026, w9027, w9028, w9029, w9030, w9031, w9032, w9033, w9034, w9035, w9036, w9037, w9038, w9039, w9040, w9041, w9042, w9043, w9044, w9045, w9046, w9047, w9048, w9049, w9050, w9051, w9052, w9053, w9054, w9055, w9056, w9057, w9058, w9059, w9060, w9061, w9062, w9063, w9064, w9065, w9066, w9067, w9068, w9069, w9070, w9071, w9072, w9073, w9074, w9075, w9076, w9077, w9078, w9079, w9080, w9081, w9082, w9083, w9084, w9085, w9086, w9087, w9088, w9089, w9090, w9091, w9092, w9093, w9094, w9095, w9096, w9097, w9098, w9099, w9100, w9101, w9102, w9103, w9104, w9105, w9106, w9107, w9108, w9109, w9110, w9111, w9112, w9113, w9114, w9115, w9116, w9117, w9118, w9119, w9120, w9121, w9122, w9123, w9124, w9125, w9126, w9127, w9128, w9129, w9130, w9131, w9132, w9133, w9134, w9135, w9136, w9137, w9138, w9139, w9140, w9141, w9142, w9143, w9144, w9145, w9146, w9147, w9148, w9149, w9150, w9151, w9152, w9153, w9154, w9155, w9156, w9157, w9158, w9159, w9160, w9161, w9162, w9163, w9164, w9165, w9166, w9167, w9168, w9169, w9170, w9171, w9172, w9173, w9174, w9175, w9176, w9177, w9178, w9179, w9180, w9181, w9182, w9183, w9184, w9185, w9186, w9187, w9188, w9189, w9190, w9191, w9192, w9193, w9194, w9195, w9196, w9197, w9198, w9199, w9200, w9201, w9202, w9203, w9204, w9205, w9206, w9207, w9208, w9209, w9210, w9211, w9212, w9213, w9214, w9215, w9216, w9217, w9218, w9219, w9220, w9221, w9222, w9223, w9224, w9225, w9226, w9227, w9228, w9229, w9230, w9231, w9232, w9233, w9234, w9235, w9236, w9237, w9238, w9239, w9240, w9241, w9242, w9243, w9244, w9245, w9246, w9247, w9248, w9249, w9250, w9251, w9252, w9253, w9254, w9255, w9256, w9257, w9258, w9259, w9260, w9261, w9262, w9263, w9264, w9265, w9266, w9267, w9268, w9269, w9270, w9271, w9272, w9273, w9274, w9275, w9276, w9277, w9278, w9279, w9280, w9281, w9282, w9283, w9284, w9285, w9286, w9287, w9288, w9289, w9290, w9291, w9292, w9293, w9294, w9295, w9296, w9297, w9298, w9299, w9300, w9301, w9302, w9303, w9304, w9305, w9306, w9307, w9308, w9309, w9310, w9311, w9312, w9313, w9314, w9315, w9316, w9317, w9318, w9319, w9320, w9321, w9322, w9323, w9324, w9325, w9326, w9327, w9328, w9329, w9330, w9331, w9332, w9333, w9334, w9335, w9336, w9337, w9338, w9339, w9340, w9341, w9342, w9343, w9344, w9345, w9346, w9347, w9348, w9349, w9350, w9351, w9352, w9353, w9354, w9355, w9356, w9357, w9358, w9359, w9360, w9361, w9362, w9363, w9364, w9365, w9366, w9367, w9368, w9369, w9370, w9371, w9372, w9373, w9374, w9375, w9376, w9377, w9378, w9379, w9380, w9381, w9382, w9383, w9384, w9385, w9386, w9387, w9388, w9389, w9390, w9391, w9392, w9393, w9394, w9395, w9396, w9397, w9398, w9399, w9400, w9401, w9402, w9403, w9404, w9405, w9406, w9407, w9408, w9409, w9410, w9411, w9412, w9413, w9414, w9415, w9416, w9417, w9418, w9419, w9420, w9421, w9422, w9423, w9424, w9425, w9426, w9427, w9428, w9429, w9430, w9431, w9432, w9433, w9434, w9435, w9436, w9437, w9438, w9439, w9440, w9441, w9442, w9443, w9444, w9445, w9446, w9447, w9448, w9449, w9450, w9451, w9452, w9453, w9454, w9455, w9456, w9457, w9458, w9459, w9460, w9461, w9462, w9463, w9464, w9465, w9466, w9467, w9468, w9469, w9470, w9471, w9472, w9473, w9474, w9475, w9476, w9477, w9478, w9479, w9480, w9481, w9482, w9483, w9484, w9485, w9486, w9487, w9488, w9489, w9490, w9491, w9492, w9493, w9494, w9495, w9496, w9497, w9498, w9499, w9500, w9501, w9502, w9503, w9504, w9505, w9506, w9507, w9508, w9509, w9510, w9511, w9512, w9513, w9514, w9515, w9516, w9517, w9518, w9519, w9520, w9521, w9522, w9523, w9524, w9525, w9526, w9527, w9528, w9529, w9530, w9531, w9532, w9533, w9534, w9535, w9536, w9537, w9538, w9539, w9540, w9541, w9542, w9543, w9544, w9545, w9546, w9547, w9548, w9549, w9550, w9551, w9552, w9553, w9554, w9555, w9556, w9557, w9558, w9559, w9560, w9561, w9562, w9563, w9564, w9565, w9566, w9567, w9568, w9569, w9570, w9571, w9572, w9573, w9574, w9575, w9576, w9577, w9578, w9579, w9580, w9581, w9582, w9583, w9584, w9585, w9586, w9587, w9588, w9589, w9590, w9591, w9592, w9593, w9594, w9595, w9596, w9597, w9598, w9599, w9600, w9601, w9602, w9603, w9604, w9605, w9606, w9607, w9608, w9609, w9610, w9611, w9612, w9613, w9614, w9615, w9616, w9617, w9618, w9619, w9620, w9621, w9622, w9623, w9624, w9625, w9626, w9627, w9628, w9629, w9630, w9631, w9632, w9633, w9634, w9635, w9636, w9637, w9638, w9639, w9640, w9641, w9642, w9643, w9644, w9645, w9646, w9647, w9648, w9649, w9650, w9651, w9652, w9653, w9654, w9655, w9656, w9657, w9658, w9659, w9660, w9661, w9662, w9663, w9664, w9665, w9666, w9667, w9668, w9669, w9670, w9671, w9672, w9673, w9674, w9675, w9676, w9677, w9678, w9679, w9680, w9681, w9682, w9683, w9684, w9685, w9686, w9687, w9688, w9689, w9690, w9691, w9692, w9693, w9694, w9695, w9696, w9697, w9698, w9699, w9700, w9701, w9702, w9703, w9704, w9705, w9706, w9707, w9708, w9709, w9710, w9711, w9712, w9713, w9714, w9715, w9716, w9717, w9718, w9719, w9720, w9721, w9722, w9723, w9724, w9725, w9726, w9727, w9728, w9729, w9730, w9731, w9732, w9733, w9734, w9735, w9736, w9737, w9738, w9739, w9740, w9741, w9742, w9743, w9744, w9745, w9746, w9747, w9748, w9749, w9750, w9751, w9752, w9753, w9754, w9755, w9756, w9757, w9758, w9759, w9760, w9761, w9762, w9763, w9764, w9765, w9766, w9767, w9768, w9769, w9770, w9771, w9772, w9773, w9774, w9775, w9776, w9777, w9778, w9779, w9780, w9781, w9782, w9783, w9784, w9785, w9786, w9787, w9788, w9789, w9790, w9791, w9792, w9793, w9794, w9795, w9796, w9797, w9798, w9799, w9800, w9801, w9802, w9803, w9804, w9805, w9806, w9807, w9808, w9809, w9810, w9811, w9812, w9813, w9814, w9815, w9816, w9817, w9818, w9819, w9820, w9821, w9822, w9823, w9824, w9825, w9826, w9827, w9828, w9829, w9830, w9831, w9832, w9833, w9834, w9835, w9836, w9837, w9838, w9839, w9840, w9841, w9842, w9843, w9844, w9845, w9846, w9847, w9848, w9849, w9850, w9851, w9852, w9853, w9854, w9855, w9856, w9857, w9858, w9859, w9860, w9861, w9862, w9863, w9864, w9865, w9866, w9867, w9868, w9869, w9870, w9871, w9872, w9873, w9874, w9875, w9876, w9877, w9878, w9879, w9880, w9881, w9882, w9883, w9884, w9885, w9886, w9887, w9888, w9889, w9890, w9891, w9892, w9893, w9894, w9895, w9896, w9897, w9898, w9899, w9900, w9901, w9902, w9903, w9904, w9905, w9906, w9907, w9908, w9909, w9910, w9911, w9912, w9913, w9914, w9915, w9916, w9917, w9918, w9919, w9920, w9921, w9922, w9923, w9924, w9925, w9926, w9927, w9928, w9929, w9930, w9931, w9932, w9933, w9934, w9935, w9936, w9937, w9938, w9939, w9940, w9941, w9942, w9943, w9944, w9945, w9946, w9947, w9948, w9949, w9950, w9951, w9952, w9953, w9954, w9955, w9956, w9957, w9958, w9959, w9960, w9961, w9962, w9963, w9964, w9965, w9966, w9967, w9968, w9969, w9970, w9971, w9972, w9973, w9974, w9975, w9976, w9977, w9978, w9979, w9980, w9981, w9982, w9983, w9984, w9985, w9986, w9987, w9988, w9989, w9990, w9991, w9992, w9993, w9994, w9995, w9996, w9997, w9998, w9999, w10000, w10001, w10002, w10003, w10004, w10005, w10006, w10007, w10008, w10009, w10010, w10011, w10012, w10013, w10014, w10015, w10016, w10017, w10018, w10019, w10020, w10021, w10022, w10023, w10024, w10025, w10026, w10027, w10028, w10029, w10030, w10031, w10032, w10033, w10034, w10035, w10036, w10037, w10038, w10039, w10040, w10041, w10042, w10043, w10044, w10045, w10046, w10047, w10048, w10049, w10050, w10051, w10052, w10053, w10054, w10055, w10056, w10057, w10058, w10059, w10060, w10061, w10062, w10063, w10064, w10065, w10066, w10067, w10068, w10069, w10070, w10071, w10072, w10073, w10074, w10075, w10076, w10077, w10078, w10079, w10080, w10081, w10082, w10083, w10084, w10085, w10086, w10087, w10088, w10089, w10090, w10091, w10092, w10093, w10094, w10095, w10096, w10097, w10098, w10099, w10100, w10101, w10102, w10103, w10104, w10105, w10106, w10107, w10108, w10109, w10110, w10111, w10112, w10113, w10114, w10115, w10116, w10117, w10118, w10119, w10120, w10121, w10122, w10123, w10124, w10125, w10126, w10127, w10128, w10129, w10130, w10131, w10132, w10133, w10134, w10135, w10136, w10137, w10138, w10139, w10140, w10141, w10142, w10143, w10144, w10145, w10146, w10147, w10148, w10149, w10150, w10151, w10152, w10153, w10154, w10155, w10156, w10157, w10158, w10159, w10160, w10161, w10162, w10163, w10164, w10165, w10166, w10167, w10168, w10169, w10170, w10171, w10172, w10173, w10174, w10175, w10176, w10177, w10178, w10179, w10180, w10181, w10182, w10183, w10184, w10185, w10186, w10187, w10188, w10189, w10190, w10191, w10192, w10193, w10194, w10195, w10196, w10197, w10198, w10199, w10200, w10201, w10202, w10203, w10204, w10205, w10206, w10207, w10208, w10209, w10210, w10211, w10212, w10213, w10214, w10215, w10216, w10217, w10218, w10219, w10220, w10221, w10222, w10223, w10224, w10225, w10226, w10227, w10228, w10229, w10230, w10231, w10232, w10233, w10234, w10235, w10236, w10237, w10238, w10239, w10240, w10241, w10242, w10243, w10244, w10245, w10246, w10247, w10248, w10249, w10250, w10251, w10252, w10253, w10254, w10255, w10256, w10257, w10258, w10259, w10260, w10261, w10262, w10263, w10264, w10265, w10266, w10267, w10268, w10269, w10270, w10271, w10272, w10273, w10274, w10275, w10276, w10277, w10278, w10279, w10280, w10281, w10282, w10283, w10284, w10285, w10286, w10287, w10288, w10289, w10290, w10291, w10292, w10293, w10294, w10295, w10296, w10297, w10298, w10299, w10300, w10301, w10302, w10303, w10304, w10305, w10306, w10307, w10308, w10309, w10310, w10311, w10312, w10313, w10314, w10315, w10316, w10317, w10318, w10319, w10320, w10321, w10322, w10323, w10324, w10325, w10326, w10327, w10328, w10329, w10330, w10331, w10332, w10333, w10334, w10335, w10336, w10337, w10338, w10339, w10340, w10341, w10342, w10343, w10344, w10345, w10346, w10347, w10348, w10349, w10350, w10351, w10352, w10353, w10354, w10355, w10356, w10357, w10358, w10359, w10360, w10361, w10362, w10363, w10364, w10365, w10366, w10367, w10368, w10369, w10370, w10371, w10372, w10373, w10374, w10375, w10376, w10377, w10378, w10379, w10380, w10381, w10382, w10383, w10384, w10385, w10386, w10387, w10388, w10389, w10390, w10391, w10392, w10393, w10394, w10395, w10396, w10397, w10398, w10399, w10400, w10401, w10402, w10403, w10404, w10405, w10406, w10407, w10408, w10409, w10410, w10411, w10412, w10413, w10414, w10415, w10416, w10417, w10418, w10419, w10420, w10421, w10422, w10423, w10424, w10425, w10426, w10427, w10428, w10429, w10430, w10431, w10432, w10433, w10434, w10435, w10436, w10437, w10438, w10439, w10440, w10441, w10442, w10443, w10444, w10445, w10446, w10447, w10448, w10449, w10450, w10451, w10452, w10453, w10454, w10455, w10456, w10457, w10458, w10459, w10460, w10461, w10462, w10463, w10464, w10465, w10466, w10467, w10468, w10469, w10470, w10471, w10472, w10473, w10474, w10475, w10476, w10477, w10478, w10479, w10480, w10481, w10482, w10483, w10484, w10485, w10486, w10487, w10488, w10489, w10490, w10491, w10492, w10493, w10494, w10495, w10496, w10497, w10498, w10499, w10500, w10501, w10502, w10503, w10504, w10505, w10506, w10507, w10508, w10509, w10510, w10511, w10512, w10513, w10514, w10515, w10516, w10517, w10518, w10519, w10520, w10521, w10522, w10523, w10524, w10525, w10526, w10527, w10528, w10529, w10530, w10531, w10532, w10533, w10534, w10535, w10536, w10537, w10538, w10539, w10540, w10541, w10542, w10543, w10544, w10545, w10546, w10547, w10548, w10549, w10550, w10551, w10552, w10553, w10554, w10555, w10556, w10557, w10558, w10559, w10560, w10561, w10562, w10563, w10564, w10565, w10566, w10567, w10568, w10569, w10570, w10571, w10572, w10573, w10574, w10575, w10576, w10577, w10578, w10579, w10580, w10581, w10582, w10583, w10584, w10585, w10586, w10587, w10588, w10589, w10590, w10591, w10592, w10593, w10594, w10595, w10596, w10597, w10598, w10599, w10600, w10601, w10602, w10603, w10604, w10605, w10606, w10607, w10608, w10609, w10610, w10611, w10612, w10613, w10614, w10615, w10616, w10617, w10618, w10619, w10620, w10621, w10622, w10623, w10624, w10625, w10626, w10627, w10628, w10629, w10630, w10631, w10632, w10633, w10634, w10635, w10636, w10637, w10638, w10639, w10640, w10641, w10642, w10643, w10644, w10645, w10646, w10647, w10648, w10649, w10650, w10651, w10652, w10653, w10654, w10655, w10656, w10657, w10658, w10659, w10660, w10661, w10662, w10663, w10664, w10665, w10666, w10667, w10668, w10669, w10670, w10671, w10672, w10673, w10674, w10675, w10676, w10677, w10678, w10679, w10680, w10681, w10682, w10683, w10684, w10685, w10686, w10687, w10688, w10689, w10690, w10691, w10692, w10693, w10694, w10695, w10696, w10697, w10698, w10699, w10700, w10701, w10702, w10703, w10704, w10705, w10706, w10707, w10708, w10709, w10710, w10711, w10712, w10713, w10714, w10715, w10716, w10717, w10718, w10719, w10720, w10721, w10722, w10723, w10724, w10725, w10726, w10727, w10728, w10729, w10730, w10731, w10732, w10733, w10734, w10735, w10736, w10737, w10738, w10739, w10740, w10741, w10742, w10743, w10744, w10745, w10746, w10747, w10748, w10749, w10750, w10751, w10752, w10753, w10754, w10755, w10756, w10757, w10758, w10759, w10760, w10761, w10762, w10763, w10764, w10765, w10766, w10767, w10768, w10769, w10770, w10771, w10772, w10773, w10774, w10775, w10776, w10777, w10778, w10779, w10780, w10781, w10782, w10783, w10784, w10785, w10786, w10787, w10788, w10789, w10790, w10791, w10792, w10793, w10794, w10795, w10796, w10797, w10798, w10799, w10800, w10801, w10802, w10803, w10804, w10805, w10806, w10807, w10808, w10809, w10810, w10811, w10812, w10813, w10814, w10815, w10816, w10817, w10818, w10819, w10820, w10821, w10822, w10823, w10824, w10825, w10826, w10827, w10828, w10829, w10830, w10831, w10832, w10833, w10834, w10835, w10836, w10837, w10838, w10839, w10840, w10841, w10842, w10843, w10844, w10845, w10846, w10847, w10848, w10849, w10850, w10851, w10852, w10853, w10854, w10855, w10856, w10857, w10858, w10859, w10860, w10861, w10862, w10863, w10864, w10865, w10866, w10867, w10868, w10869, w10870, w10871, w10872, w10873, w10874, w10875, w10876, w10877, w10878, w10879, w10880, w10881, w10882, w10883, w10884, w10885, w10886, w10887, w10888, w10889, w10890, w10891, w10892, w10893, w10894, w10895, w10896, w10897, w10898, w10899, w10900, w10901, w10902, w10903, w10904, w10905, w10906, w10907, w10908, w10909, w10910, w10911, w10912, w10913, w10914, w10915, w10916, w10917, w10918, w10919, w10920, w10921, w10922, w10923, w10924, w10925, w10926, w10927, w10928, w10929, w10930, w10931, w10932, w10933, w10934, w10935, w10936, w10937, w10938, w10939, w10940, w10941, w10942, w10943, w10944, w10945, w10946, w10947, w10948, w10949, w10950, w10951, w10952, w10953, w10954, w10955, w10956, w10957, w10958, w10959, w10960, w10961, w10962, w10963, w10964, w10965, w10966, w10967, w10968, w10969, w10970, w10971, w10972, w10973, w10974, w10975, w10976, w10977, w10978, w10979, w10980, w10981, w10982, w10983, w10984, w10985, w10986, w10987, w10988, w10989, w10990, w10991, w10992, w10993, w10994, w10995, w10996, w10997, w10998, w10999, w11000, w11001, w11002, w11003, w11004, w11005, w11006, w11007, w11008, w11009, w11010, w11011, w11012, w11013, w11014, w11015, w11016, w11017, w11018, w11019, w11020, w11021, w11022, w11023, w11024, w11025, w11026, w11027, w11028, w11029, w11030, w11031, w11032, w11033, w11034, w11035, w11036, w11037, w11038, w11039, w11040, w11041, w11042, w11043, w11044, w11045, w11046, w11047, w11048, w11049, w11050, w11051, w11052, w11053, w11054, w11055, w11056, w11057, w11058, w11059, w11060, w11061, w11062, w11063, w11064, w11065, w11066, w11067, w11068, w11069, w11070, w11071, w11072, w11073, w11074, w11075, w11076, w11077, w11078, w11079, w11080, w11081, w11082, w11083, w11084, w11085, w11086, w11087, w11088, w11089, w11090, w11091, w11092, w11093, w11094, w11095, w11096, w11097, w11098, w11099, w11100, w11101, w11102, w11103, w11104, w11105, w11106, w11107, w11108, w11109, w11110, w11111, w11112, w11113, w11114, w11115, w11116, w11117, w11118, w11119, w11120, w11121, w11122, w11123, w11124, w11125, w11126, w11127, w11128, w11129, w11130, w11131, w11132, w11133, w11134, w11135, w11136, w11137, w11138, w11139, w11140, w11141, w11142, w11143, w11144, w11145, w11146, w11147, w11148, w11149, w11150, w11151, w11152, w11153, w11154, w11155, w11156, w11157, w11158, w11159, w11160, w11161, w11162, w11163, w11164, w11165, w11166, w11167, w11168, w11169, w11170, w11171, w11172, w11173, w11174, w11175, w11176, w11177, w11178, w11179, w11180, w11181, w11182, w11183, w11184, w11185, w11186, w11187, w11188, w11189, w11190, w11191, w11192, w11193, w11194, w11195, w11196, w11197, w11198, w11199, w11200, w11201, w11202, w11203, w11204, w11205, w11206, w11207, w11208, w11209, w11210, w11211, w11212, w11213, w11214, w11215, w11216, w11217, w11218, w11219, w11220, w11221, w11222, w11223, w11224, w11225, w11226, w11227, w11228, w11229, w11230, w11231, w11232, w11233, w11234, w11235, w11236, w11237, w11238, w11239, w11240, w11241, w11242, w11243, w11244, w11245, w11246, w11247, w11248, w11249, w11250, w11251, w11252, w11253, w11254, w11255, w11256, w11257, w11258, w11259, w11260, w11261, w11262, w11263, w11264, w11265, w11266, w11267, w11268, w11269, w11270, w11271, w11272, w11273, w11274, w11275, w11276, w11277, w11278, w11279, w11280, w11281, w11282, w11283, w11284, w11285, w11286, w11287, w11288, w11289, w11290, w11291, w11292, w11293, w11294, w11295, w11296, w11297, w11298, w11299, w11300, w11301, w11302, w11303, w11304, w11305, w11306, w11307, w11308, w11309, w11310, w11311, w11312, w11313, w11314, w11315, w11316, w11317, w11318, w11319, w11320, w11321, w11322, w11323, w11324, w11325, w11326, w11327, w11328, w11329, w11330, w11331, w11332, w11333, w11334, w11335, w11336, w11337, w11338, w11339, w11340, w11341, w11342, w11343, w11344, w11345, w11346, w11347, w11348, w11349, w11350, w11351, w11352, w11353, w11354, w11355, w11356, w11357, w11358, w11359, w11360, w11361, w11362, w11363, w11364, w11365, w11366, w11367, w11368, w11369, w11370, w11371, w11372, w11373, w11374, w11375, w11376, w11377, w11378, w11379, w11380, w11381, w11382, w11383, w11384, w11385, w11386, w11387, w11388, w11389, w11390, w11391, w11392, w11393, w11394, w11395, w11396, w11397, w11398, w11399, w11400, w11401, w11402, w11403, w11404, w11405, w11406, w11407, w11408, w11409, w11410, w11411, w11412, w11413, w11414, w11415, w11416, w11417, w11418, w11419, w11420, w11421, w11422, w11423, w11424, w11425, w11426, w11427, w11428, w11429, w11430, w11431, w11432, w11433, w11434, w11435, w11436, w11437, w11438, w11439, w11440, w11441, w11442, w11443, w11444, w11445, w11446, w11447, w11448, w11449, w11450, w11451, w11452, w11453, w11454, w11455, w11456, w11457, w11458, w11459, w11460, w11461, w11462, w11463, w11464, w11465, w11466, w11467, w11468, w11469, w11470, w11471, w11472, w11473, w11474, w11475, w11476, w11477, w11478, w11479, w11480, w11481, w11482, w11483, w11484, w11485, w11486, w11487, w11488, w11489, w11490, w11491, w11492, w11493, w11494, w11495, w11496, w11497, w11498, w11499, w11500, w11501, w11502, w11503, w11504, w11505, w11506, w11507, w11508, w11509, w11510, w11511, w11512, w11513, w11514, w11515, w11516, w11517, w11518, w11519, w11520, w11521, w11522, w11523, w11524, w11525, w11526, w11527, w11528, w11529, w11530, w11531, w11532, w11533, w11534, w11535, w11536, w11537, w11538, w11539, w11540, w11541, w11542, w11543, w11544, w11545, w11546, w11547, w11548, w11549, w11550, w11551, w11552, w11553, w11554, w11555, w11556, w11557, w11558, w11559, w11560, w11561, w11562, w11563, w11564, w11565, w11566, w11567, w11568, w11569, w11570, w11571, w11572, w11573, w11574, w11575, w11576, w11577, w11578, w11579, w11580, w11581, w11582, w11583, w11584, w11585, w11586, w11587, w11588, w11589, w11590, w11591, w11592, w11593, w11594, w11595, w11596, w11597, w11598, w11599, w11600, w11601, w11602, w11603, w11604, w11605, w11606, w11607, w11608, w11609, w11610, w11611, w11612, w11613, w11614, w11615, w11616, w11617, w11618, w11619, w11620, w11621, w11622, w11623, w11624, w11625, w11626, w11627, w11628, w11629, w11630, w11631, w11632, w11633, w11634, w11635, w11636, w11637, w11638, w11639, w11640, w11641, w11642, w11643, w11644, w11645, w11646, w11647, w11648, w11649, w11650, w11651, w11652, w11653, w11654, w11655, w11656, w11657, w11658, w11659, w11660, w11661, w11662, w11663, w11664, w11665, w11666, w11667, w11668, w11669, w11670, w11671, w11672, w11673, w11674, w11675, w11676, w11677, w11678, w11679, w11680, w11681, w11682, w11683, w11684, w11685, w11686, w11687, w11688, w11689, w11690, w11691, w11692, w11693, w11694, w11695, w11696, w11697, w11698, w11699, w11700, w11701, w11702, w11703, w11704, w11705, w11706, w11707, w11708, w11709, w11710, w11711, w11712, w11713, w11714, w11715, w11716, w11717, w11718, w11719, w11720, w11721, w11722, w11723, w11724, w11725, w11726, w11727, w11728, w11729, w11730, w11731, w11732, w11733, w11734, w11735, w11736, w11737, w11738, w11739, w11740, w11741, w11742, w11743, w11744, w11745, w11746, w11747, w11748, w11749, w11750, w11751, w11752, w11753, w11754, w11755, w11756, w11757, w11758, w11759, w11760, w11761, w11762, w11763, w11764, w11765, w11766, w11767, w11768, w11769, w11770, w11771, w11772, w11773, w11774, w11775, w11776, w11777, w11778, w11779, w11780, w11781, w11782, w11783, w11784, w11785, w11786, w11787, w11788, w11789, w11790, w11791, w11792, w11793, w11794, w11795, w11796, w11797, w11798, w11799, w11800, w11801, w11802, w11803, w11804, w11805, w11806, w11807, w11808, w11809, w11810, w11811, w11812, w11813, w11814, w11815, w11816, w11817, w11818, w11819, w11820, w11821, w11822, w11823, w11824, w11825, w11826, w11827, w11828, w11829, w11830, w11831, w11832, w11833, w11834, w11835, w11836, w11837, w11838, w11839, w11840, w11841, w11842, w11843, w11844, w11845, w11846, w11847, w11848, w11849, w11850, w11851, w11852, w11853, w11854, w11855, w11856, w11857, w11858, w11859, w11860, w11861, w11862, w11863, w11864, w11865, w11866, w11867, w11868, w11869, w11870, w11871, w11872, w11873, w11874, w11875, w11876, w11877, w11878, w11879, w11880, w11881, w11882, w11883, w11884, w11885, w11886, w11887, w11888, w11889, w11890, w11891, w11892, w11893, w11894, w11895, w11896, w11897, w11898, w11899, w11900, w11901, w11902, w11903, w11904, w11905, w11906, w11907, w11908, w11909, w11910, w11911, w11912, w11913, w11914, w11915, w11916, w11917, w11918, w11919, w11920, w11921, w11922, w11923, w11924, w11925, w11926, w11927, w11928, w11929, w11930, w11931, w11932, w11933, w11934, w11935, w11936, w11937, w11938, w11939, w11940, w11941, w11942, w11943, w11944, w11945, w11946, w11947, w11948, w11949, w11950, w11951, w11952, w11953, w11954, w11955, w11956, w11957, w11958, w11959, w11960, w11961, w11962, w11963, w11964, w11965, w11966, w11967, w11968, w11969, w11970, w11971, w11972, w11973, w11974, w11975, w11976, w11977, w11978, w11979, w11980, w11981, w11982, w11983, w11984, w11985, w11986, w11987, w11988, w11989, w11990, w11991, w11992, w11993, w11994, w11995, w11996, w11997, w11998, w11999, w12000, w12001, w12002, w12003, w12004, w12005, w12006, w12007, w12008, w12009, w12010, w12011, w12012, w12013, w12014, w12015, w12016, w12017, w12018, w12019, w12020, w12021, w12022, w12023, w12024, w12025, w12026, w12027, w12028, w12029, w12030, w12031, w12032, w12033, w12034, w12035, w12036, w12037, w12038, w12039, w12040, w12041, w12042, w12043, w12044, w12045, w12046, w12047, w12048, w12049, w12050, w12051, w12052, w12053, w12054, w12055, w12056, w12057, w12058, w12059, w12060, w12061, w12062, w12063, w12064, w12065, w12066, w12067, w12068, w12069, w12070, w12071, w12072, w12073, w12074, w12075, w12076, w12077, w12078, w12079, w12080, w12081, w12082, w12083, w12084, w12085, w12086, w12087, w12088, w12089, w12090, w12091, w12092, w12093, w12094, w12095, w12096, w12097, w12098, w12099, w12100, w12101, w12102, w12103, w12104, w12105, w12106, w12107, w12108, w12109, w12110, w12111, w12112, w12113, w12114, w12115, w12116, w12117, w12118, w12119, w12120, w12121, w12122, w12123, w12124, w12125, w12126, w12127, w12128, w12129, w12130, w12131, w12132, w12133, w12134, w12135, w12136, w12137, w12138, w12139, w12140, w12141, w12142, w12143, w12144, w12145, w12146, w12147, w12148, w12149, w12150, w12151, w12152, w12153, w12154, w12155, w12156, w12157, w12158, w12159, w12160, w12161, w12162, w12163, w12164, w12165, w12166, w12167, w12168, w12169, w12170, w12171, w12172, w12173, w12174, w12175, w12176, w12177, w12178, w12179, w12180, w12181, w12182, w12183, w12184, w12185, w12186, w12187, w12188, w12189, w12190, w12191, w12192, w12193, w12194, w12195, w12196, w12197, w12198, w12199, w12200, w12201, w12202, w12203, w12204, w12205, w12206, w12207, w12208, w12209, w12210, w12211, w12212, w12213, w12214, w12215, w12216, w12217, w12218, w12219, w12220, w12221, w12222, w12223, w12224, w12225, w12226, w12227, w12228, w12229, w12230, w12231, w12232, w12233, w12234, w12235, w12236, w12237, w12238, w12239, w12240, w12241, w12242, w12243, w12244, w12245, w12246, w12247, w12248, w12249, w12250, w12251, w12252, w12253, w12254, w12255, w12256, w12257, w12258, w12259, w12260, w12261, w12262, w12263, w12264, w12265, w12266, w12267, w12268, w12269, w12270, w12271, w12272, w12273, w12274, w12275, w12276, w12277, w12278, w12279, w12280, w12281, w12282, w12283, w12284, w12285, w12286, w12287, w12288, w12289, w12290, w12291, w12292, w12293, w12294, w12295, w12296, w12297, w12298, w12299, w12300, w12301, w12302, w12303, w12304, w12305, w12306, w12307, w12308, w12309, w12310, w12311, w12312, w12313, w12314, w12315, w12316, w12317, w12318, w12319, w12320, w12321, w12322, w12323, w12324, w12325, w12326, w12327, w12328, w12329, w12330, w12331, w12332, w12333, w12334, w12335, w12336, w12337, w12338, w12339, w12340, w12341, w12342, w12343, w12344, w12345, w12346, w12347, w12348, w12349, w12350, w12351, w12352, w12353, w12354, w12355, w12356, w12357, w12358, w12359, w12360, w12361, w12362, w12363, w12364, w12365, w12366, w12367, w12368, w12369, w12370, w12371, w12372, w12373, w12374, w12375, w12376, w12377, w12378, w12379, w12380, w12381, w12382, w12383, w12384, w12385, w12386, w12387, w12388, w12389, w12390, w12391, w12392, w12393, w12394, w12395, w12396, w12397, w12398, w12399, w12400, w12401, w12402, w12403, w12404, w12405, w12406, w12407, w12408, w12409, w12410, w12411, w12412, w12413, w12414, w12415, w12416, w12417, w12418, w12419, w12420, w12421, w12422, w12423, w12424, w12425, w12426, w12427, w12428, w12429, w12430, w12431, w12432, w12433, w12434, w12435, w12436, w12437, w12438, w12439, w12440, w12441, w12442, w12443, w12444, w12445, w12446, w12447, w12448, w12449, w12450, w12451, w12452, w12453, w12454, w12455, w12456, w12457, w12458, w12459, w12460, w12461, w12462, w12463, w12464, w12465, w12466, w12467, w12468, w12469, w12470, w12471, w12472, w12473, w12474, w12475, w12476, w12477, w12478, w12479, w12480, w12481, w12482, w12483, w12484, w12485, w12486, w12487, w12488, w12489, w12490, w12491, w12492, w12493, w12494, w12495, w12496, w12497, w12498, w12499, w12500, w12501, w12502, w12503, w12504, w12505, w12506, w12507, w12508, w12509, w12510, w12511, w12512, w12513, w12514, w12515, w12516, w12517, w12518, w12519, w12520, w12521, w12522, w12523, w12524, w12525, w12526, w12527, w12528, w12529, w12530, w12531, w12532, w12533, w12534, w12535, w12536, w12537, w12538, w12539, w12540, w12541, w12542, w12543, w12544, w12545, w12546, w12547, w12548, w12549, w12550, w12551, w12552, w12553, w12554, w12555, w12556, w12557, w12558, w12559, w12560, w12561, w12562, w12563, w12564, w12565, w12566, w12567, w12568, w12569, w12570, w12571, w12572, w12573, w12574, w12575, w12576, w12577, w12578, w12579, w12580, w12581, w12582, w12583, w12584, w12585, w12586, w12587, w12588, w12589, w12590, w12591, w12592, w12593, w12594, w12595, w12596, w12597, w12598, w12599, w12600, w12601, w12602, w12603, w12604, w12605, w12606, w12607, w12608, w12609, w12610, w12611, w12612, w12613, w12614, w12615, w12616, w12617, w12618, w12619, w12620, w12621, w12622, w12623, w12624, w12625, w12626, w12627, w12628, w12629, w12630, w12631, w12632, w12633, w12634, w12635, w12636, w12637, w12638, w12639, w12640, w12641, w12642, w12643, w12644, w12645, w12646, w12647, w12648, w12649, w12650, w12651, w12652, w12653, w12654, w12655, w12656, w12657, w12658, w12659, w12660, w12661, w12662, w12663, w12664, w12665, w12666, w12667, w12668, w12669, w12670, w12671, w12672, w12673, w12674, w12675, w12676, w12677, w12678, w12679, w12680, w12681, w12682, w12683, w12684, w12685, w12686, w12687, w12688, w12689, w12690, w12691, w12692, w12693, w12694, w12695, w12696, w12697, w12698, w12699, w12700, w12701, w12702, w12703, w12704, w12705, w12706, w12707, w12708, w12709, w12710, w12711, w12712, w12713, w12714, w12715, w12716, w12717, w12718, w12719, w12720, w12721, w12722, w12723, w12724, w12725, w12726, w12727, w12728, w12729, w12730, w12731, w12732, w12733, w12734, w12735, w12736, w12737, w12738, w12739, w12740, w12741, w12742, w12743, w12744, w12745, w12746, w12747, w12748, w12749, w12750, w12751, w12752, w12753, w12754, w12755, w12756, w12757, w12758, w12759, w12760, w12761, w12762, w12763, w12764, w12765, w12766, w12767, w12768, w12769, w12770, w12771, w12772, w12773, w12774, w12775, w12776, w12777, w12778, w12779, w12780, w12781, w12782, w12783, w12784, w12785, w12786, w12787, w12788, w12789, w12790, w12791, w12792, w12793, w12794, w12795, w12796, w12797, w12798, w12799, w12800, w12801, w12802, w12803, w12804, w12805, w12806, w12807, w12808, w12809, w12810, w12811, w12812, w12813, w12814, w12815, w12816, w12817, w12818, w12819, w12820, w12821, w12822, w12823, w12824, w12825, w12826, w12827, w12828, w12829, w12830, w12831, w12832, w12833, w12834, w12835, w12836, w12837, w12838, w12839, w12840, w12841, w12842, w12843, w12844, w12845, w12846, w12847, w12848, w12849, w12850, w12851, w12852, w12853, w12854, w12855, w12856, w12857, w12858, w12859, w12860, w12861, w12862, w12863, w12864, w12865, w12866, w12867, w12868, w12869, w12870, w12871, w12872, w12873, w12874, w12875, w12876, w12877, w12878, w12879, w12880, w12881, w12882, w12883, w12884, w12885, w12886, w12887, w12888, w12889, w12890, w12891, w12892, w12893, w12894, w12895, w12896, w12897, w12898, w12899, w12900, w12901, w12902, w12903, w12904, w12905, w12906, w12907, w12908, w12909, w12910, w12911, w12912, w12913, w12914, w12915, w12916, w12917, w12918, w12919, w12920, w12921, w12922, w12923, w12924, w12925, w12926, w12927, w12928, w12929, w12930, w12931, w12932, w12933, w12934, w12935, w12936, w12937, w12938, w12939, w12940, w12941, w12942, w12943, w12944, w12945, w12946, w12947, w12948, w12949, w12950, w12951, w12952, w12953, w12954, w12955, w12956, w12957, w12958, w12959, w12960, w12961, w12962, w12963, w12964, w12965, w12966, w12967, w12968, w12969, w12970, w12971, w12972, w12973, w12974, w12975, w12976, w12977, w12978, w12979, w12980, w12981, w12982, w12983, w12984, w12985, w12986, w12987, w12988, w12989, w12990, w12991, w12992, w12993, w12994, w12995, w12996, w12997, w12998, w12999, w13000, w13001, w13002, w13003, w13004, w13005, w13006, w13007, w13008, w13009, w13010, w13011, w13012, w13013, w13014, w13015, w13016, w13017, w13018, w13019, w13020, w13021, w13022, w13023, w13024, w13025, w13026, w13027, w13028, w13029, w13030, w13031, w13032, w13033, w13034, w13035, w13036, w13037, w13038, w13039, w13040, w13041, w13042, w13043, w13044, w13045, w13046, w13047, w13048, w13049, w13050, w13051, w13052, w13053, w13054, w13055, w13056, w13057, w13058, w13059, w13060, w13061, w13062, w13063, w13064, w13065, w13066, w13067, w13068, w13069, w13070, w13071, w13072, w13073, w13074, w13075, w13076, w13077, w13078, w13079, w13080, w13081, w13082, w13083, w13084, w13085, w13086, w13087, w13088, w13089, w13090, w13091, w13092, w13093, w13094, w13095, w13096, w13097, w13098, w13099, w13100, w13101, w13102, w13103, w13104, w13105, w13106, w13107, w13108, w13109, w13110, w13111, w13112, w13113, w13114, w13115, w13116, w13117, w13118, w13119, w13120, w13121, w13122, w13123, w13124, w13125, w13126, w13127, w13128, w13129, w13130, w13131, w13132, w13133, w13134, w13135, w13136, w13137, w13138, w13139, w13140, w13141, w13142, w13143, w13144, w13145, w13146, w13147, w13148, w13149, w13150, w13151, w13152, w13153, w13154, w13155, w13156, w13157, w13158, w13159, w13160, w13161, w13162, w13163, w13164, w13165, w13166, w13167, w13168, w13169, w13170, w13171, w13172, w13173, w13174, w13175, w13176, w13177, w13178, w13179, w13180, w13181, w13182, w13183, w13184, w13185, w13186, w13187, w13188, w13189, w13190, w13191, w13192, w13193, w13194, w13195, w13196, w13197, w13198, w13199, w13200, w13201, w13202, w13203, w13204, w13205, w13206, w13207, w13208, w13209, w13210, w13211, w13212, w13213, w13214, w13215, w13216, w13217, w13218, w13219, w13220, w13221, w13222, w13223, w13224, w13225, w13226, w13227, w13228, w13229, w13230, w13231, w13232, w13233, w13234, w13235, w13236, w13237, w13238, w13239, w13240, w13241, w13242, w13243, w13244, w13245, w13246, w13247, w13248, w13249, w13250, w13251, w13252, w13253, w13254, w13255, w13256, w13257, w13258, w13259, w13260, w13261, w13262, w13263, w13264, w13265, w13266, w13267, w13268, w13269, w13270, w13271, w13272, w13273, w13274, w13275, w13276, w13277, w13278, w13279, w13280, w13281, w13282, w13283, w13284, w13285, w13286, w13287, w13288, w13289, w13290, w13291, w13292, w13293, w13294, w13295, w13296, w13297, w13298, w13299, w13300, w13301, w13302, w13303, w13304, w13305, w13306, w13307, w13308, w13309, w13310, w13311, w13312, w13313, w13314, w13315, w13316, w13317, w13318, w13319, w13320, w13321, w13322, w13323, w13324, w13325, w13326, w13327, w13328, w13329, w13330, w13331, w13332, w13333, w13334, w13335, w13336, w13337, w13338, w13339, w13340, w13341, w13342, w13343, w13344, w13345, w13346, w13347, w13348, w13349, w13350, w13351, w13352, w13353, w13354, w13355, w13356, w13357, w13358, w13359, w13360, w13361, w13362, w13363, w13364, w13365, w13366, w13367, w13368, w13369, w13370, w13371, w13372, w13373, w13374, w13375, w13376, w13377, w13378, w13379, w13380, w13381, w13382, w13383, w13384, w13385, w13386, w13387, w13388, w13389, w13390, w13391, w13392, w13393, w13394, w13395, w13396, w13397, w13398, w13399, w13400, w13401, w13402, w13403, w13404, w13405, w13406, w13407, w13408, w13409, w13410, w13411, w13412, w13413, w13414, w13415, w13416, w13417, w13418, w13419, w13420, w13421, w13422, w13423, w13424, w13425, w13426, w13427, w13428, w13429, w13430, w13431, w13432, w13433, w13434, w13435, w13436, w13437, w13438, w13439, w13440, w13441, w13442, w13443, w13444, w13445, w13446, w13447, w13448, w13449, w13450, w13451, w13452, w13453, w13454, w13455, w13456, w13457, w13458, w13459, w13460, w13461, w13462, w13463, w13464, w13465, w13466, w13467, w13468, w13469, w13470, w13471, w13472, w13473, w13474, w13475, w13476, w13477, w13478, w13479, w13480, w13481, w13482, w13483, w13484, w13485, w13486, w13487, w13488, w13489, w13490, w13491, w13492, w13493, w13494, w13495, w13496, w13497, w13498, w13499, w13500, w13501, w13502, w13503, w13504, w13505, w13506, w13507, w13508, w13509, w13510, w13511, w13512, w13513, w13514, w13515, w13516, w13517, w13518, w13519, w13520, w13521, w13522, w13523, w13524, w13525, w13526, w13527, w13528, w13529, w13530, w13531, w13532, w13533, w13534, w13535, w13536, w13537, w13538, w13539, w13540, w13541, w13542, w13543, w13544, w13545, w13546, w13547, w13548, w13549, w13550, w13551, w13552, w13553, w13554, w13555, w13556, w13557, w13558, w13559, w13560, w13561, w13562, w13563, w13564, w13565, w13566, w13567, w13568, w13569, w13570, w13571, w13572, w13573, w13574, w13575, w13576, w13577, w13578, w13579, w13580, w13581, w13582, w13583, w13584, w13585, w13586, w13587, w13588, w13589, w13590, w13591, w13592, w13593, w13594, w13595, w13596, w13597, w13598, w13599, w13600, w13601, w13602, w13603, w13604, w13605, w13606, w13607, w13608, w13609, w13610, w13611, w13612, w13613, w13614, w13615, w13616, w13617, w13618, w13619, w13620, w13621, w13622, w13623, w13624, w13625, w13626, w13627, w13628, w13629, w13630, w13631, w13632, w13633, w13634, w13635, w13636, w13637, w13638, w13639, w13640, w13641, w13642, w13643, w13644, w13645, w13646, w13647, w13648, w13649, w13650, w13651, w13652, w13653, w13654, w13655, w13656, w13657, w13658, w13659, w13660, w13661, w13662, w13663, w13664, w13665, w13666, w13667, w13668, w13669, w13670, w13671, w13672, w13673, w13674, w13675, w13676, w13677, w13678, w13679, w13680, w13681, w13682, w13683, w13684, w13685, w13686, w13687, w13688, w13689, w13690, w13691, w13692, w13693, w13694, w13695, w13696, w13697, w13698, w13699, w13700, w13701, w13702, w13703, w13704, w13705, w13706, w13707, w13708, w13709, w13710, w13711, w13712, w13713, w13714, w13715, w13716, w13717, w13718, w13719, w13720, w13721, w13722, w13723, w13724, w13725, w13726, w13727, w13728, w13729, w13730, w13731, w13732, w13733, w13734, w13735, w13736, w13737, w13738, w13739, w13740, w13741, w13742, w13743, w13744, w13745, w13746, w13747, w13748, w13749, w13750, w13751, w13752, w13753, w13754, w13755, w13756, w13757, w13758, w13759, w13760, w13761, w13762, w13763, w13764, w13765, w13766, w13767, w13768, w13769, w13770, w13771, w13772, w13773, w13774, w13775, w13776, w13777, w13778, w13779, w13780, w13781, w13782, w13783, w13784, w13785, w13786, w13787, w13788, w13789, w13790, w13791, w13792, w13793, w13794, w13795, w13796, w13797, w13798, w13799, w13800, w13801, w13802, w13803, w13804, w13805, w13806, w13807, w13808, w13809, w13810, w13811, w13812, w13813, w13814, w13815, w13816, w13817, w13818, w13819, w13820, w13821, w13822, w13823, w13824, w13825, w13826, w13827, w13828, w13829, w13830, w13831, w13832, w13833, w13834, w13835, w13836, w13837, w13838, w13839, w13840, w13841, w13842, w13843, w13844, w13845, w13846, w13847, w13848, w13849, w13850, w13851, w13852, w13853, w13854, w13855, w13856, w13857, w13858, w13859, w13860, w13861, w13862, w13863, w13864, w13865, w13866, w13867, w13868, w13869, w13870, w13871, w13872, w13873, w13874, w13875, w13876, w13877, w13878, w13879, w13880, w13881, w13882, w13883, w13884, w13885, w13886, w13887, w13888, w13889, w13890, w13891, w13892, w13893, w13894, w13895, w13896, w13897, w13898, w13899, w13900, w13901, w13902, w13903, w13904, w13905, w13906, w13907, w13908, w13909, w13910, w13911, w13912, w13913, w13914, w13915, w13916, w13917, w13918, w13919, w13920, w13921, w13922, w13923, w13924, w13925, w13926, w13927, w13928, w13929, w13930, w13931, w13932, w13933, w13934, w13935, w13936, w13937, w13938, w13939, w13940, w13941, w13942, w13943, w13944, w13945, w13946, w13947, w13948, w13949, w13950, w13951, w13952, w13953, w13954, w13955, w13956, w13957, w13958, w13959, w13960, w13961, w13962, w13963, w13964, w13965, w13966, w13967, w13968, w13969, w13970, w13971, w13972, w13973, w13974, w13975, w13976, w13977, w13978, w13979, w13980, w13981, w13982, w13983, w13984, w13985, w13986, w13987, w13988, w13989, w13990, w13991, w13992, w13993, w13994, w13995, w13996, w13997, w13998, w13999, w14000, w14001, w14002, w14003, w14004, w14005, w14006, w14007, w14008, w14009, w14010, w14011, w14012, w14013, w14014, w14015, w14016, w14017, w14018, w14019, w14020, w14021, w14022, w14023, w14024, w14025, w14026, w14027, w14028, w14029, w14030, w14031, w14032, w14033, w14034, w14035, w14036, w14037, w14038, w14039, w14040, w14041, w14042, w14043, w14044, w14045, w14046, w14047, w14048, w14049, w14050, w14051, w14052, w14053, w14054, w14055, w14056, w14057, w14058, w14059, w14060, w14061, w14062, w14063, w14064, w14065, w14066, w14067, w14068, w14069, w14070, w14071, w14072, w14073, w14074, w14075, w14076, w14077;
assign w0 = A_718 & A_719;
assign w1 = A_718 & ~A_719;
assign w2 = ~A_718 & A_719;
assign w3 = ~w1 & ~w2;
assign w4 = (~w0 & w3) | (~w0 & w13183) | (w3 & w13183);
assign w5 = A_715 & A_716;
assign w6 = A_715 & ~A_716;
assign w7 = ~A_715 & A_716;
assign w8 = ~w6 & ~w7;
assign w9 = (~w5 & w8) | (~w5 & w13184) | (w8 & w13184);
assign w10 = w4 & ~w9;
assign w11 = ~w4 & w9;
assign w12 = A_717 & ~w6;
assign w13 = ~w7 & w12;
assign w14 = ~A_717 & ~w8;
assign w15 = ~w13 & ~w14;
assign w16 = A_720 & ~w1;
assign w17 = ~w2 & w16;
assign w18 = ~A_720 & ~w3;
assign w19 = ~w17 & ~w18;
assign w20 = ~w15 & ~w19;
assign w21 = w20 & w22;
assign w22 = ~w10 & ~w11;
assign w23 = ~w20 & ~w22;
assign w24 = ~w21 & ~w23;
assign w25 = ~w15 & w19;
assign w26 = w15 & ~w19;
assign w27 = ~w25 & ~w26;
assign w28 = w20 & ~w22;
assign w29 = ~w4 & ~w9;
assign w30 = ~w28 & ~w29;
assign w31 = ~w27 & ~w30;
assign w32 = ~w24 & ~w31;
assign w33 = ~w24 & ~w30;
assign w34 = A_724 & A_725;
assign w35 = A_724 & ~A_725;
assign w36 = ~A_724 & A_725;
assign w37 = ~w35 & ~w36;
assign w38 = (~w34 & w37) | (~w34 & w13185) | (w37 & w13185);
assign w39 = A_721 & A_722;
assign w40 = A_721 & ~A_722;
assign w41 = ~A_721 & A_722;
assign w42 = ~w40 & ~w41;
assign w43 = (~w39 & w42) | (~w39 & w13186) | (w42 & w13186);
assign w44 = ~w38 & w43;
assign w45 = w38 & ~w43;
assign w46 = ~w44 & ~w45;
assign w47 = A_723 & ~w40;
assign w48 = ~w41 & w47;
assign w49 = ~A_723 & ~w42;
assign w50 = ~w48 & ~w49;
assign w51 = A_726 & ~w35;
assign w52 = ~w36 & w51;
assign w53 = ~A_726 & ~w37;
assign w54 = ~w52 & ~w53;
assign w55 = ~w50 & ~w54;
assign w56 = ~w46 & w55;
assign w57 = ~w38 & ~w43;
assign w58 = ~w56 & ~w57;
assign w59 = w55 & w46;
assign w60 = ~w46 & ~w55;
assign w61 = ~w59 & ~w60;
assign w62 = ~w58 & ~w61;
assign w63 = ~w50 & w54;
assign w64 = w50 & ~w54;
assign w65 = ~w63 & ~w64;
assign w66 = ~w27 & ~w65;
assign w67 = ~w62 & w66;
assign w68 = ~w33 & w67;
assign w69 = ~w58 & ~w65;
assign w70 = ~w61 & ~w69;
assign w71 = ~w68 & ~w70;
assign w72 = ~w61 & w66;
assign w73 = ~w62 & w72;
assign w74 = ~w33 & ~w69;
assign w75 = w73 & w74;
assign w76 = (w32 & w71) | (w32 & w13653) | (w71 & w13653);
assign w77 = ~w68 & w70;
assign w78 = w68 & ~w70;
assign w79 = ~w77 & ~w78;
assign w80 = ~w32 & ~w79;
assign w81 = ~w62 & ~w65;
assign w82 = ~w27 & ~w33;
assign w83 = ~w81 & w82;
assign w84 = w81 & ~w82;
assign w85 = ~w83 & ~w84;
assign w86 = ~A_709 & A_710;
assign w87 = A_709 & ~A_710;
assign w88 = A_711 & ~w87;
assign w89 = ~w86 & w88;
assign w90 = ~w86 & ~w87;
assign w91 = ~A_711 & ~w90;
assign w92 = ~w89 & ~w91;
assign w93 = ~A_712 & A_713;
assign w94 = A_712 & ~A_713;
assign w95 = A_714 & ~w94;
assign w96 = ~w93 & w95;
assign w97 = ~w93 & ~w94;
assign w98 = ~A_714 & ~w97;
assign w99 = ~w96 & ~w98;
assign w100 = ~w92 & w99;
assign w101 = w92 & ~w99;
assign w102 = ~w100 & ~w101;
assign w103 = A_712 & A_713;
assign w104 = (~w103 & w97) | (~w103 & w13187) | (w97 & w13187);
assign w105 = A_709 & A_710;
assign w106 = (~w105 & w90) | (~w105 & w13188) | (w90 & w13188);
assign w107 = ~w104 & w106;
assign w108 = w104 & ~w106;
assign w109 = ~w107 & ~w108;
assign w110 = ~w92 & ~w99;
assign w111 = ~w109 & w110;
assign w112 = ~w104 & ~w106;
assign w113 = ~w111 & ~w112;
assign w114 = w110 & w109;
assign w115 = ~w109 & ~w110;
assign w116 = ~w114 & ~w115;
assign w117 = ~w113 & ~w116;
assign w118 = ~w102 & ~w117;
assign w119 = ~A_703 & A_704;
assign w120 = A_703 & ~A_704;
assign w121 = A_705 & ~w120;
assign w122 = ~w119 & w121;
assign w123 = ~w119 & ~w120;
assign w124 = ~A_705 & ~w123;
assign w125 = ~w122 & ~w124;
assign w126 = ~A_706 & A_707;
assign w127 = A_706 & ~A_707;
assign w128 = A_708 & ~w127;
assign w129 = ~w126 & w128;
assign w130 = ~w126 & ~w127;
assign w131 = ~A_708 & ~w130;
assign w132 = ~w129 & ~w131;
assign w133 = ~w125 & w132;
assign w134 = w125 & ~w132;
assign w135 = ~w133 & ~w134;
assign w136 = A_706 & A_707;
assign w137 = (~w136 & w130) | (~w136 & w13189) | (w130 & w13189);
assign w138 = A_703 & A_704;
assign w139 = (~w138 & w123) | (~w138 & w13190) | (w123 & w13190);
assign w140 = ~w137 & w139;
assign w141 = w137 & ~w139;
assign w142 = ~w140 & ~w141;
assign w143 = ~w125 & ~w132;
assign w144 = ~w142 & w143;
assign w145 = ~w137 & ~w139;
assign w146 = ~w144 & ~w145;
assign w147 = w143 & w142;
assign w148 = ~w142 & ~w143;
assign w149 = ~w147 & ~w148;
assign w150 = ~w146 & ~w149;
assign w151 = ~w135 & ~w150;
assign w152 = ~w118 & w151;
assign w153 = w118 & ~w151;
assign w154 = ~w152 & ~w153;
assign w155 = ~w85 & ~w154;
assign w156 = ~w80 & w13654;
assign w157 = (~w155 & w80) | (~w155 & w13655) | (w80 & w13655);
assign w158 = ~w156 & ~w157;
assign w159 = ~w135 & ~w146;
assign w160 = ~w149 & ~w159;
assign w161 = ~w102 & ~w135;
assign w162 = ~w117 & w161;
assign w163 = ~w150 & w162;
assign w164 = ~w102 & ~w113;
assign w165 = ~w116 & ~w164;
assign w166 = ~w163 & w165;
assign w167 = w163 & ~w165;
assign w168 = ~w166 & ~w167;
assign w169 = ~w160 & ~w168;
assign w170 = ~w163 & ~w165;
assign w171 = ~w116 & w161;
assign w172 = ~w117 & w171;
assign w173 = ~w150 & ~w164;
assign w174 = w172 & w173;
assign w175 = (w160 & w170) | (w160 & w13797) | (w170 & w13797);
assign w176 = ~w169 & ~w175;
assign w177 = ~w158 & w176;
assign w178 = ~w80 & w13656;
assign w179 = (w155 & w80) | (w155 & w13798) | (w80 & w13798);
assign w180 = (~w176 & w179) | (~w176 & w13657) | (w179 & w13657);
assign w181 = ~w177 & ~w180;
assign w182 = A_730 & A_731;
assign w183 = A_730 & ~A_731;
assign w184 = ~A_730 & A_731;
assign w185 = ~w183 & ~w184;
assign w186 = (~w182 & w185) | (~w182 & w13191) | (w185 & w13191);
assign w187 = A_727 & A_728;
assign w188 = A_727 & ~A_728;
assign w189 = ~A_727 & A_728;
assign w190 = ~w188 & ~w189;
assign w191 = (~w187 & w190) | (~w187 & w13192) | (w190 & w13192);
assign w192 = w186 & ~w191;
assign w193 = ~w186 & w191;
assign w194 = A_729 & ~w188;
assign w195 = ~w189 & w194;
assign w196 = ~A_729 & ~w190;
assign w197 = ~w195 & ~w196;
assign w198 = A_732 & ~w183;
assign w199 = ~w184 & w198;
assign w200 = ~A_732 & ~w185;
assign w201 = ~w199 & ~w200;
assign w202 = ~w197 & ~w201;
assign w203 = w202 & w204;
assign w204 = ~w192 & ~w193;
assign w205 = ~w202 & ~w204;
assign w206 = ~w203 & ~w205;
assign w207 = ~w197 & w201;
assign w208 = w197 & ~w201;
assign w209 = ~w207 & ~w208;
assign w210 = w202 & ~w204;
assign w211 = ~w186 & ~w191;
assign w212 = ~w210 & ~w211;
assign w213 = ~w209 & ~w212;
assign w214 = ~w206 & ~w213;
assign w215 = ~w206 & ~w212;
assign w216 = A_736 & A_737;
assign w217 = A_736 & ~A_737;
assign w218 = ~A_736 & A_737;
assign w219 = ~w217 & ~w218;
assign w220 = (~w216 & w219) | (~w216 & w13193) | (w219 & w13193);
assign w221 = A_733 & A_734;
assign w222 = A_733 & ~A_734;
assign w223 = ~A_733 & A_734;
assign w224 = ~w222 & ~w223;
assign w225 = (~w221 & w224) | (~w221 & w13194) | (w224 & w13194);
assign w226 = ~w220 & w225;
assign w227 = w220 & ~w225;
assign w228 = ~w226 & ~w227;
assign w229 = A_735 & ~w222;
assign w230 = ~w223 & w229;
assign w231 = ~A_735 & ~w224;
assign w232 = ~w230 & ~w231;
assign w233 = A_738 & ~w217;
assign w234 = ~w218 & w233;
assign w235 = ~A_738 & ~w219;
assign w236 = ~w234 & ~w235;
assign w237 = ~w232 & ~w236;
assign w238 = ~w228 & w237;
assign w239 = ~w220 & ~w225;
assign w240 = ~w238 & ~w239;
assign w241 = w237 & w228;
assign w242 = ~w228 & ~w237;
assign w243 = ~w241 & ~w242;
assign w244 = ~w240 & ~w243;
assign w245 = ~w232 & w236;
assign w246 = w232 & ~w236;
assign w247 = ~w245 & ~w246;
assign w248 = ~w209 & ~w247;
assign w249 = ~w244 & w248;
assign w250 = ~w215 & w249;
assign w251 = ~w240 & ~w247;
assign w252 = ~w243 & ~w251;
assign w253 = ~w250 & w252;
assign w254 = w250 & ~w252;
assign w255 = ~w253 & ~w254;
assign w256 = ~w214 & ~w255;
assign w257 = ~w250 & ~w252;
assign w258 = ~w243 & w248;
assign w259 = ~w244 & w258;
assign w260 = ~w215 & ~w251;
assign w261 = w259 & w260;
assign w262 = (w214 & w257) | (w214 & w13658) | (w257 & w13658);
assign w263 = ~w256 & ~w262;
assign w264 = A_742 & A_743;
assign w265 = A_742 & ~A_743;
assign w266 = ~A_742 & A_743;
assign w267 = ~w265 & ~w266;
assign w268 = (~w264 & w267) | (~w264 & w13195) | (w267 & w13195);
assign w269 = A_739 & A_740;
assign w270 = A_739 & ~A_740;
assign w271 = ~A_739 & A_740;
assign w272 = ~w270 & ~w271;
assign w273 = (~w269 & w272) | (~w269 & w13196) | (w272 & w13196);
assign w274 = w268 & ~w273;
assign w275 = ~w268 & w273;
assign w276 = A_741 & ~w270;
assign w277 = ~w271 & w276;
assign w278 = ~A_741 & ~w272;
assign w279 = ~w277 & ~w278;
assign w280 = A_744 & ~w265;
assign w281 = ~w266 & w280;
assign w282 = ~A_744 & ~w267;
assign w283 = ~w281 & ~w282;
assign w284 = ~w279 & ~w283;
assign w285 = w284 & w286;
assign w286 = ~w274 & ~w275;
assign w287 = ~w284 & ~w286;
assign w288 = ~w285 & ~w287;
assign w289 = ~w279 & w283;
assign w290 = w279 & ~w283;
assign w291 = ~w289 & ~w290;
assign w292 = w284 & ~w286;
assign w293 = ~w268 & ~w273;
assign w294 = ~w292 & ~w293;
assign w295 = ~w291 & ~w294;
assign w296 = ~w288 & ~w295;
assign w297 = ~w288 & ~w294;
assign w298 = A_748 & A_749;
assign w299 = A_748 & ~A_749;
assign w300 = ~A_748 & A_749;
assign w301 = ~w299 & ~w300;
assign w302 = (~w298 & w301) | (~w298 & w13197) | (w301 & w13197);
assign w303 = A_745 & A_746;
assign w304 = A_745 & ~A_746;
assign w305 = ~A_745 & A_746;
assign w306 = ~w304 & ~w305;
assign w307 = (~w303 & w306) | (~w303 & w13198) | (w306 & w13198);
assign w308 = ~w302 & w307;
assign w309 = w302 & ~w307;
assign w310 = ~w308 & ~w309;
assign w311 = A_747 & ~w304;
assign w312 = ~w305 & w311;
assign w313 = ~A_747 & ~w306;
assign w314 = ~w312 & ~w313;
assign w315 = A_750 & ~w299;
assign w316 = ~w300 & w315;
assign w317 = ~A_750 & ~w301;
assign w318 = ~w316 & ~w317;
assign w319 = ~w314 & ~w318;
assign w320 = ~w310 & w319;
assign w321 = ~w302 & ~w307;
assign w322 = ~w320 & ~w321;
assign w323 = w319 & w310;
assign w324 = ~w310 & ~w319;
assign w325 = ~w323 & ~w324;
assign w326 = ~w322 & ~w325;
assign w327 = ~w314 & w318;
assign w328 = w314 & ~w318;
assign w329 = ~w327 & ~w328;
assign w330 = ~w291 & ~w329;
assign w331 = ~w326 & w330;
assign w332 = ~w297 & w331;
assign w333 = ~w322 & ~w329;
assign w334 = ~w325 & ~w333;
assign w335 = ~w332 & ~w334;
assign w336 = ~w325 & w330;
assign w337 = ~w326 & w336;
assign w338 = ~w297 & ~w333;
assign w339 = w337 & w338;
assign w340 = (w296 & w335) | (w296 & w13478) | (w335 & w13478);
assign w341 = ~w332 & w334;
assign w342 = w332 & ~w334;
assign w343 = ~w341 & ~w342;
assign w344 = ~w296 & ~w343;
assign w345 = ~w326 & ~w329;
assign w346 = ~w291 & ~w297;
assign w347 = ~w345 & w346;
assign w348 = w345 & ~w346;
assign w349 = ~w347 & ~w348;
assign w350 = ~w244 & ~w247;
assign w351 = ~w209 & ~w215;
assign w352 = ~w350 & w351;
assign w353 = w350 & ~w351;
assign w354 = ~w352 & ~w353;
assign w355 = ~w349 & ~w354;
assign w356 = ~w344 & w13479;
assign w357 = (w355 & w344) | (w355 & w13480) | (w344 & w13480);
assign w358 = ~w356 & ~w357;
assign w359 = ~w263 & ~w358;
assign w360 = ~w344 & w13481;
assign w361 = (~w355 & w344) | (~w355 & w13659) | (w344 & w13659);
assign w362 = (w263 & w361) | (w263 & w13482) | (w361 & w13482);
assign w363 = ~w349 & w354;
assign w364 = w349 & ~w354;
assign w365 = ~w363 & ~w364;
assign w366 = ~w85 & w154;
assign w367 = w85 & ~w154;
assign w368 = ~w366 & ~w367;
assign w369 = ~w365 & ~w368;
assign w370 = ~w369 & ~w362;
assign w371 = ~w359 & w370;
assign w372 = ~w359 & ~w362;
assign w373 = w369 & ~w372;
assign w374 = (~w181 & w373) | (~w181 & w13799) | (w373 & w13799);
assign w375 = w369 & ~w362;
assign w376 = ~w359 & w375;
assign w377 = ~w369 & ~w372;
assign w378 = (w181 & w377) | (w181 & w13660) | (w377 & w13660);
assign w379 = ~w365 & w368;
assign w380 = w365 & ~w368;
assign w381 = ~w379 & ~w380;
assign w382 = ~A_697 & A_698;
assign w383 = A_697 & ~A_698;
assign w384 = A_699 & ~w383;
assign w385 = ~w382 & w384;
assign w386 = ~w382 & ~w383;
assign w387 = ~A_699 & ~w386;
assign w388 = ~w385 & ~w387;
assign w389 = ~A_700 & A_701;
assign w390 = A_700 & ~A_701;
assign w391 = A_702 & ~w390;
assign w392 = ~w389 & w391;
assign w393 = ~w389 & ~w390;
assign w394 = ~A_702 & ~w393;
assign w395 = ~w392 & ~w394;
assign w396 = ~w388 & w395;
assign w397 = w388 & ~w395;
assign w398 = ~w396 & ~w397;
assign w399 = A_700 & A_701;
assign w400 = (~w399 & w393) | (~w399 & w13199) | (w393 & w13199);
assign w401 = A_697 & A_698;
assign w402 = (~w401 & w386) | (~w401 & w13200) | (w386 & w13200);
assign w403 = ~w400 & w402;
assign w404 = w400 & ~w402;
assign w405 = ~w403 & ~w404;
assign w406 = ~w388 & ~w395;
assign w407 = ~w405 & w406;
assign w408 = ~w400 & ~w402;
assign w409 = ~w407 & ~w408;
assign w410 = w406 & w405;
assign w411 = ~w405 & ~w406;
assign w412 = ~w410 & ~w411;
assign w413 = ~w409 & ~w412;
assign w414 = ~w398 & ~w413;
assign w415 = ~A_691 & A_692;
assign w416 = A_691 & ~A_692;
assign w417 = A_693 & ~w416;
assign w418 = ~w415 & w417;
assign w419 = ~w415 & ~w416;
assign w420 = ~A_693 & ~w419;
assign w421 = ~w418 & ~w420;
assign w422 = ~A_694 & A_695;
assign w423 = A_694 & ~A_695;
assign w424 = A_696 & ~w423;
assign w425 = ~w422 & w424;
assign w426 = ~w422 & ~w423;
assign w427 = ~A_696 & ~w426;
assign w428 = ~w425 & ~w427;
assign w429 = ~w421 & w428;
assign w430 = w421 & ~w428;
assign w431 = ~w429 & ~w430;
assign w432 = A_694 & A_695;
assign w433 = (~w432 & w426) | (~w432 & w13201) | (w426 & w13201);
assign w434 = A_691 & A_692;
assign w435 = (~w434 & w419) | (~w434 & w13202) | (w419 & w13202);
assign w436 = ~w433 & w435;
assign w437 = w433 & ~w435;
assign w438 = ~w436 & ~w437;
assign w439 = ~w421 & ~w428;
assign w440 = ~w438 & w439;
assign w441 = ~w433 & ~w435;
assign w442 = ~w440 & ~w441;
assign w443 = w439 & w438;
assign w444 = ~w438 & ~w439;
assign w445 = ~w443 & ~w444;
assign w446 = ~w442 & ~w445;
assign w447 = ~w431 & ~w446;
assign w448 = ~w414 & w447;
assign w449 = w414 & ~w447;
assign w450 = ~w448 & ~w449;
assign w451 = ~A_685 & A_686;
assign w452 = A_685 & ~A_686;
assign w453 = A_687 & ~w452;
assign w454 = ~w451 & w453;
assign w455 = ~w451 & ~w452;
assign w456 = ~A_687 & ~w455;
assign w457 = ~w454 & ~w456;
assign w458 = ~A_688 & A_689;
assign w459 = A_688 & ~A_689;
assign w460 = A_690 & ~w459;
assign w461 = ~w458 & w460;
assign w462 = ~w458 & ~w459;
assign w463 = ~A_690 & ~w462;
assign w464 = ~w461 & ~w463;
assign w465 = ~w457 & w464;
assign w466 = w457 & ~w464;
assign w467 = ~w465 & ~w466;
assign w468 = A_688 & A_689;
assign w469 = (~w468 & w462) | (~w468 & w13203) | (w462 & w13203);
assign w470 = A_685 & A_686;
assign w471 = (~w470 & w455) | (~w470 & w13204) | (w455 & w13204);
assign w472 = ~w469 & w471;
assign w473 = w469 & ~w471;
assign w474 = ~w472 & ~w473;
assign w475 = ~w457 & ~w464;
assign w476 = ~w474 & w475;
assign w477 = ~w469 & ~w471;
assign w478 = ~w476 & ~w477;
assign w479 = w475 & w474;
assign w480 = ~w474 & ~w475;
assign w481 = ~w479 & ~w480;
assign w482 = ~w478 & ~w481;
assign w483 = ~w467 & ~w482;
assign w484 = ~A_679 & A_680;
assign w485 = A_679 & ~A_680;
assign w486 = A_681 & ~w485;
assign w487 = ~w484 & w486;
assign w488 = ~w484 & ~w485;
assign w489 = ~A_681 & ~w488;
assign w490 = ~w487 & ~w489;
assign w491 = ~A_682 & A_683;
assign w492 = A_682 & ~A_683;
assign w493 = A_684 & ~w492;
assign w494 = ~w491 & w493;
assign w495 = ~w491 & ~w492;
assign w496 = ~A_684 & ~w495;
assign w497 = ~w494 & ~w496;
assign w498 = ~w490 & w497;
assign w499 = w490 & ~w497;
assign w500 = ~w498 & ~w499;
assign w501 = A_682 & A_683;
assign w502 = (~w501 & w495) | (~w501 & w13205) | (w495 & w13205);
assign w503 = A_679 & A_680;
assign w504 = (~w503 & w488) | (~w503 & w13206) | (w488 & w13206);
assign w505 = ~w502 & w504;
assign w506 = w502 & ~w504;
assign w507 = ~w505 & ~w506;
assign w508 = ~w490 & ~w497;
assign w509 = ~w507 & w508;
assign w510 = ~w502 & ~w504;
assign w511 = ~w509 & ~w510;
assign w512 = w508 & w507;
assign w513 = ~w507 & ~w508;
assign w514 = ~w512 & ~w513;
assign w515 = ~w511 & ~w514;
assign w516 = ~w500 & ~w515;
assign w517 = ~w483 & w516;
assign w518 = w483 & ~w516;
assign w519 = ~w517 & ~w518;
assign w520 = ~w450 & w519;
assign w521 = w450 & ~w519;
assign w522 = ~w520 & ~w521;
assign w523 = ~A_673 & A_674;
assign w524 = A_673 & ~A_674;
assign w525 = A_675 & ~w524;
assign w526 = ~w523 & w525;
assign w527 = ~w523 & ~w524;
assign w528 = ~A_675 & ~w527;
assign w529 = ~w526 & ~w528;
assign w530 = ~A_676 & A_677;
assign w531 = A_676 & ~A_677;
assign w532 = A_678 & ~w531;
assign w533 = ~w530 & w532;
assign w534 = ~w530 & ~w531;
assign w535 = ~A_678 & ~w534;
assign w536 = ~w533 & ~w535;
assign w537 = ~w529 & w536;
assign w538 = w529 & ~w536;
assign w539 = ~w537 & ~w538;
assign w540 = A_676 & A_677;
assign w541 = (~w540 & w534) | (~w540 & w13207) | (w534 & w13207);
assign w542 = A_673 & A_674;
assign w543 = (~w542 & w527) | (~w542 & w13208) | (w527 & w13208);
assign w544 = ~w541 & w543;
assign w545 = w541 & ~w543;
assign w546 = ~w544 & ~w545;
assign w547 = ~w529 & ~w536;
assign w548 = ~w546 & w547;
assign w549 = ~w541 & ~w543;
assign w550 = ~w548 & ~w549;
assign w551 = w547 & w546;
assign w552 = ~w546 & ~w547;
assign w553 = ~w551 & ~w552;
assign w554 = ~w550 & ~w553;
assign w555 = ~w539 & ~w554;
assign w556 = ~A_667 & A_668;
assign w557 = A_667 & ~A_668;
assign w558 = A_669 & ~w557;
assign w559 = ~w556 & w558;
assign w560 = ~w556 & ~w557;
assign w561 = ~A_669 & ~w560;
assign w562 = ~w559 & ~w561;
assign w563 = ~A_670 & A_671;
assign w564 = A_670 & ~A_671;
assign w565 = A_672 & ~w564;
assign w566 = ~w563 & w565;
assign w567 = ~w563 & ~w564;
assign w568 = ~A_672 & ~w567;
assign w569 = ~w566 & ~w568;
assign w570 = ~w562 & w569;
assign w571 = w562 & ~w569;
assign w572 = ~w570 & ~w571;
assign w573 = A_670 & A_671;
assign w574 = (~w573 & w567) | (~w573 & w13209) | (w567 & w13209);
assign w575 = A_667 & A_668;
assign w576 = (~w575 & w560) | (~w575 & w13210) | (w560 & w13210);
assign w577 = ~w574 & w576;
assign w578 = w574 & ~w576;
assign w579 = ~w577 & ~w578;
assign w580 = ~w562 & ~w569;
assign w581 = ~w579 & w580;
assign w582 = ~w574 & ~w576;
assign w583 = ~w581 & ~w582;
assign w584 = w580 & w579;
assign w585 = ~w579 & ~w580;
assign w586 = ~w584 & ~w585;
assign w587 = ~w583 & ~w586;
assign w588 = ~w572 & ~w587;
assign w589 = ~w555 & w588;
assign w590 = w555 & ~w588;
assign w591 = ~w589 & ~w590;
assign w592 = ~A_661 & A_662;
assign w593 = A_661 & ~A_662;
assign w594 = A_663 & ~w593;
assign w595 = ~w592 & w594;
assign w596 = ~w592 & ~w593;
assign w597 = ~A_663 & ~w596;
assign w598 = ~w595 & ~w597;
assign w599 = ~A_664 & A_665;
assign w600 = A_664 & ~A_665;
assign w601 = A_666 & ~w600;
assign w602 = ~w599 & w601;
assign w603 = ~w599 & ~w600;
assign w604 = ~A_666 & ~w603;
assign w605 = ~w602 & ~w604;
assign w606 = ~w598 & w605;
assign w607 = w598 & ~w605;
assign w608 = ~w606 & ~w607;
assign w609 = A_664 & A_665;
assign w610 = (~w609 & w603) | (~w609 & w13211) | (w603 & w13211);
assign w611 = A_661 & A_662;
assign w612 = (~w611 & w596) | (~w611 & w13212) | (w596 & w13212);
assign w613 = ~w610 & w612;
assign w614 = w610 & ~w612;
assign w615 = ~w613 & ~w614;
assign w616 = ~w598 & ~w605;
assign w617 = ~w615 & w616;
assign w618 = ~w610 & ~w612;
assign w619 = ~w617 & ~w618;
assign w620 = w616 & w615;
assign w621 = ~w615 & ~w616;
assign w622 = ~w620 & ~w621;
assign w623 = ~w619 & ~w622;
assign w624 = ~w608 & ~w623;
assign w625 = ~A_655 & A_656;
assign w626 = A_655 & ~A_656;
assign w627 = A_657 & ~w626;
assign w628 = ~w625 & w627;
assign w629 = ~w625 & ~w626;
assign w630 = ~A_657 & ~w629;
assign w631 = ~w628 & ~w630;
assign w632 = ~A_658 & A_659;
assign w633 = A_658 & ~A_659;
assign w634 = A_660 & ~w633;
assign w635 = ~w632 & w634;
assign w636 = ~w632 & ~w633;
assign w637 = ~A_660 & ~w636;
assign w638 = ~w635 & ~w637;
assign w639 = ~w631 & w638;
assign w640 = w631 & ~w638;
assign w641 = ~w639 & ~w640;
assign w642 = A_658 & A_659;
assign w643 = (~w642 & w636) | (~w642 & w13213) | (w636 & w13213);
assign w644 = A_655 & A_656;
assign w645 = (~w644 & w629) | (~w644 & w13214) | (w629 & w13214);
assign w646 = ~w643 & w645;
assign w647 = w643 & ~w645;
assign w648 = ~w646 & ~w647;
assign w649 = ~w631 & ~w638;
assign w650 = ~w648 & w649;
assign w651 = ~w643 & ~w645;
assign w652 = ~w650 & ~w651;
assign w653 = w649 & w648;
assign w654 = ~w648 & ~w649;
assign w655 = ~w653 & ~w654;
assign w656 = ~w652 & ~w655;
assign w657 = ~w641 & ~w656;
assign w658 = ~w624 & w657;
assign w659 = w624 & ~w657;
assign w660 = ~w658 & ~w659;
assign w661 = ~w591 & w660;
assign w662 = w591 & ~w660;
assign w663 = ~w661 & ~w662;
assign w664 = ~w522 & w663;
assign w665 = w522 & ~w663;
assign w666 = ~w664 & ~w665;
assign w667 = ~w381 & ~w666;
assign w668 = ~w378 & w667;
assign w669 = ~w374 & w668;
assign w670 = ~w374 & ~w378;
assign w671 = ~w667 & ~w670;
assign w672 = ~w669 & ~w671;
assign w673 = ~w500 & ~w511;
assign w674 = ~w514 & ~w673;
assign w675 = ~w467 & ~w500;
assign w676 = ~w482 & w675;
assign w677 = ~w515 & w676;
assign w678 = ~w467 & ~w478;
assign w679 = ~w481 & ~w678;
assign w680 = ~w677 & w679;
assign w681 = w677 & ~w679;
assign w682 = ~w680 & ~w681;
assign w683 = ~w674 & ~w682;
assign w684 = ~w677 & ~w679;
assign w685 = ~w481 & w675;
assign w686 = ~w482 & w685;
assign w687 = ~w515 & ~w678;
assign w688 = w686 & w687;
assign w689 = (w674 & w684) | (w674 & w13661) | (w684 & w13661);
assign w690 = ~w683 & ~w689;
assign w691 = ~w431 & ~w442;
assign w692 = ~w445 & ~w691;
assign w693 = ~w398 & ~w431;
assign w694 = ~w413 & w693;
assign w695 = ~w446 & w694;
assign w696 = ~w398 & ~w409;
assign w697 = ~w412 & ~w696;
assign w698 = ~w695 & ~w697;
assign w699 = ~w412 & w693;
assign w700 = ~w413 & w699;
assign w701 = ~w446 & ~w696;
assign w702 = w700 & w701;
assign w703 = (w692 & w698) | (w692 & w13483) | (w698 & w13483);
assign w704 = ~w695 & w697;
assign w705 = w695 & ~w697;
assign w706 = ~w704 & ~w705;
assign w707 = ~w692 & ~w706;
assign w708 = ~w450 & ~w519;
assign w709 = ~w707 & w13484;
assign w710 = (w708 & w707) | (w708 & w13662) | (w707 & w13662);
assign w711 = ~w709 & ~w710;
assign w712 = ~w690 & ~w711;
assign w713 = ~w707 & w13485;
assign w714 = (~w708 & w707) | (~w708 & w13663) | (w707 & w13663);
assign w715 = (w690 & w714) | (w690 & w13486) | (w714 & w13486);
assign w716 = ~w522 & ~w663;
assign w717 = w716 & ~w715;
assign w718 = ~w712 & w717;
assign w719 = ~w712 & ~w715;
assign w720 = ~w716 & ~w719;
assign w721 = ~w572 & ~w583;
assign w722 = ~w586 & ~w721;
assign w723 = ~w539 & ~w572;
assign w724 = ~w554 & w723;
assign w725 = ~w587 & w724;
assign w726 = ~w539 & ~w550;
assign w727 = ~w553 & ~w726;
assign w728 = ~w725 & ~w727;
assign w729 = ~w553 & w723;
assign w730 = ~w554 & w729;
assign w731 = ~w587 & ~w726;
assign w732 = w730 & w731;
assign w733 = (w722 & w728) | (w722 & w13664) | (w728 & w13664);
assign w734 = ~w725 & w727;
assign w735 = w725 & ~w727;
assign w736 = ~w734 & ~w735;
assign w737 = ~w722 & ~w736;
assign w738 = ~w591 & ~w660;
assign w739 = ~w737 & w13665;
assign w740 = (~w738 & w737) | (~w738 & w13666) | (w737 & w13666);
assign w741 = ~w739 & ~w740;
assign w742 = ~w641 & ~w652;
assign w743 = ~w655 & ~w742;
assign w744 = ~w608 & ~w641;
assign w745 = ~w623 & w744;
assign w746 = ~w656 & w745;
assign w747 = ~w608 & ~w619;
assign w748 = ~w622 & ~w747;
assign w749 = ~w746 & w748;
assign w750 = w746 & ~w748;
assign w751 = ~w749 & ~w750;
assign w752 = ~w743 & ~w751;
assign w753 = ~w746 & ~w748;
assign w754 = ~w622 & w744;
assign w755 = ~w623 & w754;
assign w756 = ~w656 & ~w747;
assign w757 = w755 & w756;
assign w758 = (w743 & w753) | (w743 & w13800) | (w753 & w13800);
assign w759 = ~w752 & ~w758;
assign w760 = ~w741 & w759;
assign w761 = ~w737 & w13667;
assign w762 = (w738 & w737) | (w738 & w13801) | (w737 & w13801);
assign w763 = (~w759 & w762) | (~w759 & w13668) | (w762 & w13668);
assign w764 = ~w760 & ~w763;
assign w765 = (w764 & w720) | (w764 & w13802) | (w720 & w13802);
assign w766 = ~w716 & ~w715;
assign w767 = ~w712 & w766;
assign w768 = w716 & ~w719;
assign w769 = (~w764 & w768) | (~w764 & w13803) | (w768 & w13803);
assign w770 = ~w765 & ~w769;
assign w771 = ~w672 & w770;
assign w772 = ~w378 & ~w667;
assign w773 = ~w374 & w772;
assign w774 = w667 & ~w670;
assign w775 = ~w773 & ~w774;
assign w776 = ~w770 & ~w775;
assign w777 = ~w771 & ~w776;
assign w778 = A_778 & A_779;
assign w779 = A_778 & ~A_779;
assign w780 = ~A_778 & A_779;
assign w781 = ~w779 & ~w780;
assign w782 = (~w778 & w781) | (~w778 & w13215) | (w781 & w13215);
assign w783 = A_775 & A_776;
assign w784 = A_775 & ~A_776;
assign w785 = ~A_775 & A_776;
assign w786 = ~w784 & ~w785;
assign w787 = (~w783 & w786) | (~w783 & w13216) | (w786 & w13216);
assign w788 = w782 & ~w787;
assign w789 = ~w782 & w787;
assign w790 = A_777 & ~w784;
assign w791 = ~w785 & w790;
assign w792 = ~A_777 & ~w786;
assign w793 = ~w791 & ~w792;
assign w794 = A_780 & ~w779;
assign w795 = ~w780 & w794;
assign w796 = ~A_780 & ~w781;
assign w797 = ~w795 & ~w796;
assign w798 = ~w793 & ~w797;
assign w799 = w798 & w800;
assign w800 = ~w788 & ~w789;
assign w801 = ~w798 & ~w800;
assign w802 = ~w799 & ~w801;
assign w803 = ~w793 & w797;
assign w804 = w793 & ~w797;
assign w805 = ~w803 & ~w804;
assign w806 = w798 & ~w800;
assign w807 = ~w782 & ~w787;
assign w808 = ~w806 & ~w807;
assign w809 = ~w805 & ~w808;
assign w810 = ~w802 & ~w809;
assign w811 = ~w802 & ~w808;
assign w812 = A_784 & A_785;
assign w813 = A_784 & ~A_785;
assign w814 = ~A_784 & A_785;
assign w815 = ~w813 & ~w814;
assign w816 = (~w812 & w815) | (~w812 & w13217) | (w815 & w13217);
assign w817 = A_781 & A_782;
assign w818 = A_781 & ~A_782;
assign w819 = ~A_781 & A_782;
assign w820 = ~w818 & ~w819;
assign w821 = (~w817 & w820) | (~w817 & w13218) | (w820 & w13218);
assign w822 = ~w816 & w821;
assign w823 = w816 & ~w821;
assign w824 = ~w822 & ~w823;
assign w825 = A_783 & ~w818;
assign w826 = ~w819 & w825;
assign w827 = ~A_783 & ~w820;
assign w828 = ~w826 & ~w827;
assign w829 = A_786 & ~w813;
assign w830 = ~w814 & w829;
assign w831 = ~A_786 & ~w815;
assign w832 = ~w830 & ~w831;
assign w833 = ~w828 & ~w832;
assign w834 = ~w824 & w833;
assign w835 = ~w816 & ~w821;
assign w836 = ~w834 & ~w835;
assign w837 = w833 & w824;
assign w838 = ~w824 & ~w833;
assign w839 = ~w837 & ~w838;
assign w840 = ~w836 & ~w839;
assign w841 = ~w828 & w832;
assign w842 = w828 & ~w832;
assign w843 = ~w841 & ~w842;
assign w844 = ~w805 & ~w843;
assign w845 = ~w840 & w844;
assign w846 = ~w811 & w845;
assign w847 = ~w836 & ~w843;
assign w848 = ~w839 & ~w847;
assign w849 = ~w846 & w848;
assign w850 = w846 & ~w848;
assign w851 = ~w849 & ~w850;
assign w852 = ~w810 & ~w851;
assign w853 = ~w846 & ~w848;
assign w854 = ~w839 & w844;
assign w855 = ~w840 & w854;
assign w856 = ~w811 & ~w847;
assign w857 = w855 & w856;
assign w858 = (w810 & w853) | (w810 & w13669) | (w853 & w13669);
assign w859 = ~w852 & ~w858;
assign w860 = A_790 & A_791;
assign w861 = A_790 & ~A_791;
assign w862 = ~A_790 & A_791;
assign w863 = ~w861 & ~w862;
assign w864 = (~w860 & w863) | (~w860 & w13219) | (w863 & w13219);
assign w865 = A_787 & A_788;
assign w866 = A_787 & ~A_788;
assign w867 = ~A_787 & A_788;
assign w868 = ~w866 & ~w867;
assign w869 = (~w865 & w868) | (~w865 & w13220) | (w868 & w13220);
assign w870 = w864 & ~w869;
assign w871 = ~w864 & w869;
assign w872 = A_789 & ~w866;
assign w873 = ~w867 & w872;
assign w874 = ~A_789 & ~w868;
assign w875 = ~w873 & ~w874;
assign w876 = A_792 & ~w861;
assign w877 = ~w862 & w876;
assign w878 = ~A_792 & ~w863;
assign w879 = ~w877 & ~w878;
assign w880 = ~w875 & ~w879;
assign w881 = w880 & w882;
assign w882 = ~w870 & ~w871;
assign w883 = ~w880 & ~w882;
assign w884 = ~w881 & ~w883;
assign w885 = ~w875 & w879;
assign w886 = w875 & ~w879;
assign w887 = ~w885 & ~w886;
assign w888 = w880 & ~w882;
assign w889 = ~w864 & ~w869;
assign w890 = ~w888 & ~w889;
assign w891 = ~w887 & ~w890;
assign w892 = ~w884 & ~w891;
assign w893 = ~w884 & ~w890;
assign w894 = A_796 & A_797;
assign w895 = A_796 & ~A_797;
assign w896 = ~A_796 & A_797;
assign w897 = ~w895 & ~w896;
assign w898 = (~w894 & w897) | (~w894 & w13221) | (w897 & w13221);
assign w899 = A_793 & A_794;
assign w900 = A_793 & ~A_794;
assign w901 = ~A_793 & A_794;
assign w902 = ~w900 & ~w901;
assign w903 = (~w899 & w902) | (~w899 & w13222) | (w902 & w13222);
assign w904 = ~w898 & w903;
assign w905 = w898 & ~w903;
assign w906 = ~w904 & ~w905;
assign w907 = A_795 & ~w900;
assign w908 = ~w901 & w907;
assign w909 = ~A_795 & ~w902;
assign w910 = ~w908 & ~w909;
assign w911 = A_798 & ~w895;
assign w912 = ~w896 & w911;
assign w913 = ~A_798 & ~w897;
assign w914 = ~w912 & ~w913;
assign w915 = ~w910 & ~w914;
assign w916 = ~w906 & w915;
assign w917 = ~w898 & ~w903;
assign w918 = ~w916 & ~w917;
assign w919 = w915 & w906;
assign w920 = ~w906 & ~w915;
assign w921 = ~w919 & ~w920;
assign w922 = ~w918 & ~w921;
assign w923 = ~w910 & w914;
assign w924 = w910 & ~w914;
assign w925 = ~w923 & ~w924;
assign w926 = ~w887 & ~w925;
assign w927 = ~w922 & w926;
assign w928 = ~w893 & w927;
assign w929 = ~w918 & ~w925;
assign w930 = ~w921 & ~w929;
assign w931 = ~w928 & ~w930;
assign w932 = ~w921 & w926;
assign w933 = ~w922 & w932;
assign w934 = ~w893 & ~w929;
assign w935 = w933 & w934;
assign w936 = (w892 & w931) | (w892 & w13487) | (w931 & w13487);
assign w937 = ~w928 & w930;
assign w938 = w928 & ~w930;
assign w939 = ~w937 & ~w938;
assign w940 = ~w892 & ~w939;
assign w941 = ~w922 & ~w925;
assign w942 = ~w887 & ~w893;
assign w943 = ~w941 & w942;
assign w944 = w941 & ~w942;
assign w945 = ~w943 & ~w944;
assign w946 = ~w840 & ~w843;
assign w947 = ~w805 & ~w811;
assign w948 = ~w946 & w947;
assign w949 = w946 & ~w947;
assign w950 = ~w948 & ~w949;
assign w951 = ~w945 & ~w950;
assign w952 = ~w940 & w13488;
assign w953 = (w951 & w940) | (w951 & w13670) | (w940 & w13670);
assign w954 = ~w952 & ~w953;
assign w955 = ~w859 & ~w954;
assign w956 = ~w940 & w13489;
assign w957 = (~w951 & w940) | (~w951 & w13671) | (w940 & w13671);
assign w958 = (w859 & w957) | (w859 & w13490) | (w957 & w13490);
assign w959 = ~w945 & w950;
assign w960 = w945 & ~w950;
assign w961 = ~w959 & ~w960;
assign w962 = ~A_769 & A_770;
assign w963 = A_769 & ~A_770;
assign w964 = A_771 & ~w963;
assign w965 = ~w962 & w964;
assign w966 = ~w962 & ~w963;
assign w967 = ~A_771 & ~w966;
assign w968 = ~w965 & ~w967;
assign w969 = ~A_772 & A_773;
assign w970 = A_772 & ~A_773;
assign w971 = A_774 & ~w970;
assign w972 = ~w969 & w971;
assign w973 = ~w969 & ~w970;
assign w974 = ~A_774 & ~w973;
assign w975 = ~w972 & ~w974;
assign w976 = ~w968 & w975;
assign w977 = w968 & ~w975;
assign w978 = ~w976 & ~w977;
assign w979 = A_772 & A_773;
assign w980 = (~w979 & w973) | (~w979 & w13223) | (w973 & w13223);
assign w981 = A_769 & A_770;
assign w982 = (~w981 & w966) | (~w981 & w13224) | (w966 & w13224);
assign w983 = ~w980 & w982;
assign w984 = w980 & ~w982;
assign w985 = ~w983 & ~w984;
assign w986 = ~w968 & ~w975;
assign w987 = ~w985 & w986;
assign w988 = ~w980 & ~w982;
assign w989 = ~w987 & ~w988;
assign w990 = w986 & w985;
assign w991 = ~w985 & ~w986;
assign w992 = ~w990 & ~w991;
assign w993 = ~w989 & ~w992;
assign w994 = ~w978 & ~w993;
assign w995 = ~A_763 & A_764;
assign w996 = A_763 & ~A_764;
assign w997 = A_765 & ~w996;
assign w998 = ~w995 & w997;
assign w999 = ~w995 & ~w996;
assign w1000 = ~A_765 & ~w999;
assign w1001 = ~w998 & ~w1000;
assign w1002 = ~A_766 & A_767;
assign w1003 = A_766 & ~A_767;
assign w1004 = A_768 & ~w1003;
assign w1005 = ~w1002 & w1004;
assign w1006 = ~w1002 & ~w1003;
assign w1007 = ~A_768 & ~w1006;
assign w1008 = ~w1005 & ~w1007;
assign w1009 = ~w1001 & w1008;
assign w1010 = w1001 & ~w1008;
assign w1011 = ~w1009 & ~w1010;
assign w1012 = A_766 & A_767;
assign w1013 = (~w1012 & w1006) | (~w1012 & w13225) | (w1006 & w13225);
assign w1014 = A_763 & A_764;
assign w1015 = (~w1014 & w999) | (~w1014 & w13226) | (w999 & w13226);
assign w1016 = ~w1013 & w1015;
assign w1017 = w1013 & ~w1015;
assign w1018 = ~w1016 & ~w1017;
assign w1019 = ~w1001 & ~w1008;
assign w1020 = ~w1018 & w1019;
assign w1021 = ~w1013 & ~w1015;
assign w1022 = ~w1020 & ~w1021;
assign w1023 = w1019 & w1018;
assign w1024 = ~w1018 & ~w1019;
assign w1025 = ~w1023 & ~w1024;
assign w1026 = ~w1022 & ~w1025;
assign w1027 = ~w1011 & ~w1026;
assign w1028 = ~w994 & w1027;
assign w1029 = w994 & ~w1027;
assign w1030 = ~w1028 & ~w1029;
assign w1031 = ~A_757 & A_758;
assign w1032 = A_757 & ~A_758;
assign w1033 = A_759 & ~w1032;
assign w1034 = ~w1031 & w1033;
assign w1035 = ~w1031 & ~w1032;
assign w1036 = ~A_759 & ~w1035;
assign w1037 = ~w1034 & ~w1036;
assign w1038 = ~A_760 & A_761;
assign w1039 = A_760 & ~A_761;
assign w1040 = A_762 & ~w1039;
assign w1041 = ~w1038 & w1040;
assign w1042 = ~w1038 & ~w1039;
assign w1043 = ~A_762 & ~w1042;
assign w1044 = ~w1041 & ~w1043;
assign w1045 = ~w1037 & w1044;
assign w1046 = w1037 & ~w1044;
assign w1047 = ~w1045 & ~w1046;
assign w1048 = A_760 & A_761;
assign w1049 = (~w1048 & w1042) | (~w1048 & w13227) | (w1042 & w13227);
assign w1050 = A_757 & A_758;
assign w1051 = (~w1050 & w1035) | (~w1050 & w13228) | (w1035 & w13228);
assign w1052 = ~w1049 & w1051;
assign w1053 = w1049 & ~w1051;
assign w1054 = ~w1052 & ~w1053;
assign w1055 = ~w1037 & ~w1044;
assign w1056 = ~w1054 & w1055;
assign w1057 = ~w1049 & ~w1051;
assign w1058 = ~w1056 & ~w1057;
assign w1059 = w1055 & w1054;
assign w1060 = ~w1054 & ~w1055;
assign w1061 = ~w1059 & ~w1060;
assign w1062 = ~w1058 & ~w1061;
assign w1063 = ~w1047 & ~w1062;
assign w1064 = ~A_751 & A_752;
assign w1065 = A_751 & ~A_752;
assign w1066 = A_753 & ~w1065;
assign w1067 = ~w1064 & w1066;
assign w1068 = ~w1064 & ~w1065;
assign w1069 = ~A_753 & ~w1068;
assign w1070 = ~w1067 & ~w1069;
assign w1071 = ~A_754 & A_755;
assign w1072 = A_754 & ~A_755;
assign w1073 = A_756 & ~w1072;
assign w1074 = ~w1071 & w1073;
assign w1075 = ~w1071 & ~w1072;
assign w1076 = ~A_756 & ~w1075;
assign w1077 = ~w1074 & ~w1076;
assign w1078 = ~w1070 & w1077;
assign w1079 = w1070 & ~w1077;
assign w1080 = ~w1078 & ~w1079;
assign w1081 = A_754 & A_755;
assign w1082 = (~w1081 & w1075) | (~w1081 & w13229) | (w1075 & w13229);
assign w1083 = A_751 & A_752;
assign w1084 = (~w1083 & w1068) | (~w1083 & w13230) | (w1068 & w13230);
assign w1085 = ~w1082 & w1084;
assign w1086 = w1082 & ~w1084;
assign w1087 = ~w1085 & ~w1086;
assign w1088 = ~w1070 & ~w1077;
assign w1089 = ~w1087 & w1088;
assign w1090 = ~w1082 & ~w1084;
assign w1091 = ~w1089 & ~w1090;
assign w1092 = w1088 & w1087;
assign w1093 = ~w1087 & ~w1088;
assign w1094 = ~w1092 & ~w1093;
assign w1095 = ~w1091 & ~w1094;
assign w1096 = ~w1080 & ~w1095;
assign w1097 = ~w1063 & w1096;
assign w1098 = w1063 & ~w1096;
assign w1099 = ~w1097 & ~w1098;
assign w1100 = ~w1030 & w1099;
assign w1101 = w1030 & ~w1099;
assign w1102 = ~w1100 & ~w1101;
assign w1103 = ~w961 & ~w1102;
assign w1104 = w1103 & ~w958;
assign w1105 = ~w955 & w1104;
assign w1106 = ~w955 & ~w958;
assign w1107 = ~w1103 & ~w1106;
assign w1108 = ~w1011 & ~w1022;
assign w1109 = ~w1025 & ~w1108;
assign w1110 = ~w978 & ~w1011;
assign w1111 = ~w993 & w1110;
assign w1112 = ~w1026 & w1111;
assign w1113 = ~w978 & ~w989;
assign w1114 = ~w992 & ~w1113;
assign w1115 = ~w1112 & ~w1114;
assign w1116 = ~w992 & w1110;
assign w1117 = ~w993 & w1116;
assign w1118 = ~w1026 & ~w1113;
assign w1119 = w1117 & w1118;
assign w1120 = (w1109 & w1115) | (w1109 & w13672) | (w1115 & w13672);
assign w1121 = ~w1112 & w1114;
assign w1122 = w1112 & ~w1114;
assign w1123 = ~w1121 & ~w1122;
assign w1124 = ~w1109 & ~w1123;
assign w1125 = ~w1030 & ~w1099;
assign w1126 = ~w1124 & w13673;
assign w1127 = (~w1125 & w1124) | (~w1125 & w13674) | (w1124 & w13674);
assign w1128 = ~w1126 & ~w1127;
assign w1129 = ~w1080 & ~w1091;
assign w1130 = ~w1094 & ~w1129;
assign w1131 = ~w1047 & ~w1080;
assign w1132 = ~w1062 & w1131;
assign w1133 = ~w1095 & w1132;
assign w1134 = ~w1047 & ~w1058;
assign w1135 = ~w1061 & ~w1134;
assign w1136 = ~w1133 & w1135;
assign w1137 = w1133 & ~w1135;
assign w1138 = ~w1136 & ~w1137;
assign w1139 = ~w1130 & ~w1138;
assign w1140 = ~w1133 & ~w1135;
assign w1141 = ~w1061 & w1131;
assign w1142 = ~w1062 & w1141;
assign w1143 = ~w1095 & ~w1134;
assign w1144 = w1142 & w1143;
assign w1145 = (w1130 & w1140) | (w1130 & w13804) | (w1140 & w13804);
assign w1146 = ~w1139 & ~w1145;
assign w1147 = ~w1128 & w1146;
assign w1148 = ~w1124 & w13675;
assign w1149 = (w1125 & w1124) | (w1125 & w13805) | (w1124 & w13805);
assign w1150 = (~w1146 & w1149) | (~w1146 & w13676) | (w1149 & w13676);
assign w1151 = ~w1147 & ~w1150;
assign w1152 = (w1151 & w1107) | (w1151 & w13806) | (w1107 & w13806);
assign w1153 = ~w1103 & ~w958;
assign w1154 = ~w955 & w1153;
assign w1155 = w1103 & ~w1106;
assign w1156 = (~w1151 & w1155) | (~w1151 & w13807) | (w1155 & w13807);
assign w1157 = ~w1152 & ~w1156;
assign w1158 = A_814 & A_815;
assign w1159 = A_814 & ~A_815;
assign w1160 = ~A_814 & A_815;
assign w1161 = ~w1159 & ~w1160;
assign w1162 = (~w1158 & w1161) | (~w1158 & w13231) | (w1161 & w13231);
assign w1163 = A_811 & A_812;
assign w1164 = A_811 & ~A_812;
assign w1165 = ~A_811 & A_812;
assign w1166 = ~w1164 & ~w1165;
assign w1167 = (~w1163 & w1166) | (~w1163 & w13232) | (w1166 & w13232);
assign w1168 = w1162 & ~w1167;
assign w1169 = ~w1162 & w1167;
assign w1170 = A_813 & ~w1164;
assign w1171 = ~w1165 & w1170;
assign w1172 = ~A_813 & ~w1166;
assign w1173 = ~w1171 & ~w1172;
assign w1174 = A_816 & ~w1159;
assign w1175 = ~w1160 & w1174;
assign w1176 = ~A_816 & ~w1161;
assign w1177 = ~w1175 & ~w1176;
assign w1178 = ~w1173 & ~w1177;
assign w1179 = w1178 & w1180;
assign w1180 = ~w1168 & ~w1169;
assign w1181 = ~w1178 & ~w1180;
assign w1182 = ~w1179 & ~w1181;
assign w1183 = ~w1173 & w1177;
assign w1184 = w1173 & ~w1177;
assign w1185 = ~w1183 & ~w1184;
assign w1186 = w1178 & ~w1180;
assign w1187 = ~w1162 & ~w1167;
assign w1188 = ~w1186 & ~w1187;
assign w1189 = ~w1185 & ~w1188;
assign w1190 = ~w1182 & ~w1189;
assign w1191 = ~w1182 & ~w1188;
assign w1192 = A_820 & A_821;
assign w1193 = A_820 & ~A_821;
assign w1194 = ~A_820 & A_821;
assign w1195 = ~w1193 & ~w1194;
assign w1196 = (~w1192 & w1195) | (~w1192 & w13233) | (w1195 & w13233);
assign w1197 = A_817 & A_818;
assign w1198 = A_817 & ~A_818;
assign w1199 = ~A_817 & A_818;
assign w1200 = ~w1198 & ~w1199;
assign w1201 = (~w1197 & w1200) | (~w1197 & w13234) | (w1200 & w13234);
assign w1202 = ~w1196 & w1201;
assign w1203 = w1196 & ~w1201;
assign w1204 = ~w1202 & ~w1203;
assign w1205 = A_819 & ~w1198;
assign w1206 = ~w1199 & w1205;
assign w1207 = ~A_819 & ~w1200;
assign w1208 = ~w1206 & ~w1207;
assign w1209 = A_822 & ~w1193;
assign w1210 = ~w1194 & w1209;
assign w1211 = ~A_822 & ~w1195;
assign w1212 = ~w1210 & ~w1211;
assign w1213 = ~w1208 & ~w1212;
assign w1214 = ~w1204 & w1213;
assign w1215 = ~w1196 & ~w1201;
assign w1216 = ~w1214 & ~w1215;
assign w1217 = w1213 & w1204;
assign w1218 = ~w1204 & ~w1213;
assign w1219 = ~w1217 & ~w1218;
assign w1220 = ~w1216 & ~w1219;
assign w1221 = ~w1208 & w1212;
assign w1222 = w1208 & ~w1212;
assign w1223 = ~w1221 & ~w1222;
assign w1224 = ~w1185 & ~w1223;
assign w1225 = ~w1220 & w1224;
assign w1226 = ~w1191 & w1225;
assign w1227 = ~w1216 & ~w1223;
assign w1228 = ~w1219 & ~w1227;
assign w1229 = ~w1226 & ~w1228;
assign w1230 = ~w1219 & w1224;
assign w1231 = ~w1220 & w1230;
assign w1232 = ~w1191 & ~w1227;
assign w1233 = w1231 & w1232;
assign w1234 = (w1190 & w1229) | (w1190 & w13677) | (w1229 & w13677);
assign w1235 = ~w1226 & w1228;
assign w1236 = w1226 & ~w1228;
assign w1237 = ~w1235 & ~w1236;
assign w1238 = ~w1190 & ~w1237;
assign w1239 = ~w1220 & ~w1223;
assign w1240 = ~w1185 & ~w1191;
assign w1241 = ~w1239 & w1240;
assign w1242 = w1239 & ~w1240;
assign w1243 = ~w1241 & ~w1242;
assign w1244 = ~A_805 & A_806;
assign w1245 = A_805 & ~A_806;
assign w1246 = A_807 & ~w1245;
assign w1247 = ~w1244 & w1246;
assign w1248 = ~w1244 & ~w1245;
assign w1249 = ~A_807 & ~w1248;
assign w1250 = ~w1247 & ~w1249;
assign w1251 = ~A_808 & A_809;
assign w1252 = A_808 & ~A_809;
assign w1253 = A_810 & ~w1252;
assign w1254 = ~w1251 & w1253;
assign w1255 = ~w1251 & ~w1252;
assign w1256 = ~A_810 & ~w1255;
assign w1257 = ~w1254 & ~w1256;
assign w1258 = ~w1250 & w1257;
assign w1259 = w1250 & ~w1257;
assign w1260 = ~w1258 & ~w1259;
assign w1261 = A_808 & A_809;
assign w1262 = (~w1261 & w1255) | (~w1261 & w13235) | (w1255 & w13235);
assign w1263 = A_805 & A_806;
assign w1264 = (~w1263 & w1248) | (~w1263 & w13236) | (w1248 & w13236);
assign w1265 = ~w1262 & w1264;
assign w1266 = w1262 & ~w1264;
assign w1267 = ~w1265 & ~w1266;
assign w1268 = ~w1250 & ~w1257;
assign w1269 = ~w1267 & w1268;
assign w1270 = ~w1262 & ~w1264;
assign w1271 = ~w1269 & ~w1270;
assign w1272 = w1268 & w1267;
assign w1273 = ~w1267 & ~w1268;
assign w1274 = ~w1272 & ~w1273;
assign w1275 = ~w1271 & ~w1274;
assign w1276 = ~w1260 & ~w1275;
assign w1277 = ~A_799 & A_800;
assign w1278 = A_799 & ~A_800;
assign w1279 = A_801 & ~w1278;
assign w1280 = ~w1277 & w1279;
assign w1281 = ~w1277 & ~w1278;
assign w1282 = ~A_801 & ~w1281;
assign w1283 = ~w1280 & ~w1282;
assign w1284 = ~A_802 & A_803;
assign w1285 = A_802 & ~A_803;
assign w1286 = A_804 & ~w1285;
assign w1287 = ~w1284 & w1286;
assign w1288 = ~w1284 & ~w1285;
assign w1289 = ~A_804 & ~w1288;
assign w1290 = ~w1287 & ~w1289;
assign w1291 = ~w1283 & w1290;
assign w1292 = w1283 & ~w1290;
assign w1293 = ~w1291 & ~w1292;
assign w1294 = A_802 & A_803;
assign w1295 = (~w1294 & w1288) | (~w1294 & w13237) | (w1288 & w13237);
assign w1296 = A_799 & A_800;
assign w1297 = (~w1296 & w1281) | (~w1296 & w13238) | (w1281 & w13238);
assign w1298 = ~w1295 & w1297;
assign w1299 = w1295 & ~w1297;
assign w1300 = ~w1298 & ~w1299;
assign w1301 = ~w1283 & ~w1290;
assign w1302 = ~w1300 & w1301;
assign w1303 = ~w1295 & ~w1297;
assign w1304 = ~w1302 & ~w1303;
assign w1305 = w1301 & w1300;
assign w1306 = ~w1300 & ~w1301;
assign w1307 = ~w1305 & ~w1306;
assign w1308 = ~w1304 & ~w1307;
assign w1309 = ~w1293 & ~w1308;
assign w1310 = ~w1276 & w1309;
assign w1311 = w1276 & ~w1309;
assign w1312 = ~w1310 & ~w1311;
assign w1313 = ~w1243 & ~w1312;
assign w1314 = ~w1238 & w13678;
assign w1315 = (~w1313 & w1238) | (~w1313 & w13679) | (w1238 & w13679);
assign w1316 = ~w1314 & ~w1315;
assign w1317 = ~w1293 & ~w1304;
assign w1318 = ~w1307 & ~w1317;
assign w1319 = ~w1260 & ~w1293;
assign w1320 = ~w1275 & w1319;
assign w1321 = ~w1308 & w1320;
assign w1322 = ~w1260 & ~w1271;
assign w1323 = ~w1274 & ~w1322;
assign w1324 = ~w1321 & w1323;
assign w1325 = w1321 & ~w1323;
assign w1326 = ~w1324 & ~w1325;
assign w1327 = ~w1318 & ~w1326;
assign w1328 = ~w1321 & ~w1323;
assign w1329 = ~w1274 & w1319;
assign w1330 = ~w1275 & w1329;
assign w1331 = ~w1308 & ~w1322;
assign w1332 = w1330 & w1331;
assign w1333 = (w1318 & w1328) | (w1318 & w13808) | (w1328 & w13808);
assign w1334 = ~w1327 & ~w1333;
assign w1335 = ~w1316 & w1334;
assign w1336 = ~w1238 & w13680;
assign w1337 = (w1313 & w1238) | (w1313 & w13809) | (w1238 & w13809);
assign w1338 = (~w1334 & w1337) | (~w1334 & w13681) | (w1337 & w13681);
assign w1339 = ~w1335 & ~w1338;
assign w1340 = A_826 & A_827;
assign w1341 = A_826 & ~A_827;
assign w1342 = ~A_826 & A_827;
assign w1343 = ~w1341 & ~w1342;
assign w1344 = (~w1340 & w1343) | (~w1340 & w13239) | (w1343 & w13239);
assign w1345 = A_823 & A_824;
assign w1346 = A_823 & ~A_824;
assign w1347 = ~A_823 & A_824;
assign w1348 = ~w1346 & ~w1347;
assign w1349 = (~w1345 & w1348) | (~w1345 & w13240) | (w1348 & w13240);
assign w1350 = w1344 & ~w1349;
assign w1351 = ~w1344 & w1349;
assign w1352 = A_825 & ~w1346;
assign w1353 = ~w1347 & w1352;
assign w1354 = ~A_825 & ~w1348;
assign w1355 = ~w1353 & ~w1354;
assign w1356 = A_828 & ~w1341;
assign w1357 = ~w1342 & w1356;
assign w1358 = ~A_828 & ~w1343;
assign w1359 = ~w1357 & ~w1358;
assign w1360 = ~w1355 & ~w1359;
assign w1361 = w1360 & w1362;
assign w1362 = ~w1350 & ~w1351;
assign w1363 = ~w1360 & ~w1362;
assign w1364 = ~w1361 & ~w1363;
assign w1365 = ~w1355 & w1359;
assign w1366 = w1355 & ~w1359;
assign w1367 = ~w1365 & ~w1366;
assign w1368 = w1360 & ~w1362;
assign w1369 = ~w1344 & ~w1349;
assign w1370 = ~w1368 & ~w1369;
assign w1371 = ~w1367 & ~w1370;
assign w1372 = ~w1364 & ~w1371;
assign w1373 = ~w1364 & ~w1370;
assign w1374 = A_832 & A_833;
assign w1375 = A_832 & ~A_833;
assign w1376 = ~A_832 & A_833;
assign w1377 = ~w1375 & ~w1376;
assign w1378 = (~w1374 & w1377) | (~w1374 & w13241) | (w1377 & w13241);
assign w1379 = A_829 & A_830;
assign w1380 = A_829 & ~A_830;
assign w1381 = ~A_829 & A_830;
assign w1382 = ~w1380 & ~w1381;
assign w1383 = (~w1379 & w1382) | (~w1379 & w13242) | (w1382 & w13242);
assign w1384 = ~w1378 & w1383;
assign w1385 = w1378 & ~w1383;
assign w1386 = ~w1384 & ~w1385;
assign w1387 = A_831 & ~w1380;
assign w1388 = ~w1381 & w1387;
assign w1389 = ~A_831 & ~w1382;
assign w1390 = ~w1388 & ~w1389;
assign w1391 = A_834 & ~w1375;
assign w1392 = ~w1376 & w1391;
assign w1393 = ~A_834 & ~w1377;
assign w1394 = ~w1392 & ~w1393;
assign w1395 = ~w1390 & ~w1394;
assign w1396 = ~w1386 & w1395;
assign w1397 = ~w1378 & ~w1383;
assign w1398 = ~w1396 & ~w1397;
assign w1399 = w1395 & w1386;
assign w1400 = ~w1386 & ~w1395;
assign w1401 = ~w1399 & ~w1400;
assign w1402 = ~w1398 & ~w1401;
assign w1403 = ~w1390 & w1394;
assign w1404 = w1390 & ~w1394;
assign w1405 = ~w1403 & ~w1404;
assign w1406 = ~w1367 & ~w1405;
assign w1407 = ~w1402 & w1406;
assign w1408 = ~w1373 & w1407;
assign w1409 = ~w1398 & ~w1405;
assign w1410 = ~w1401 & ~w1409;
assign w1411 = ~w1408 & w1410;
assign w1412 = w1408 & ~w1410;
assign w1413 = ~w1411 & ~w1412;
assign w1414 = ~w1372 & ~w1413;
assign w1415 = ~w1408 & ~w1410;
assign w1416 = ~w1401 & w1406;
assign w1417 = ~w1402 & w1416;
assign w1418 = ~w1373 & ~w1409;
assign w1419 = w1417 & w1418;
assign w1420 = (w1372 & w1415) | (w1372 & w13682) | (w1415 & w13682);
assign w1421 = ~w1414 & ~w1420;
assign w1422 = A_838 & A_839;
assign w1423 = A_838 & ~A_839;
assign w1424 = ~A_838 & A_839;
assign w1425 = ~w1423 & ~w1424;
assign w1426 = (~w1422 & w1425) | (~w1422 & w13243) | (w1425 & w13243);
assign w1427 = A_835 & A_836;
assign w1428 = A_835 & ~A_836;
assign w1429 = ~A_835 & A_836;
assign w1430 = ~w1428 & ~w1429;
assign w1431 = (~w1427 & w1430) | (~w1427 & w13244) | (w1430 & w13244);
assign w1432 = w1426 & ~w1431;
assign w1433 = ~w1426 & w1431;
assign w1434 = A_837 & ~w1428;
assign w1435 = ~w1429 & w1434;
assign w1436 = ~A_837 & ~w1430;
assign w1437 = ~w1435 & ~w1436;
assign w1438 = A_840 & ~w1423;
assign w1439 = ~w1424 & w1438;
assign w1440 = ~A_840 & ~w1425;
assign w1441 = ~w1439 & ~w1440;
assign w1442 = ~w1437 & ~w1441;
assign w1443 = w1442 & w1444;
assign w1444 = ~w1432 & ~w1433;
assign w1445 = ~w1442 & ~w1444;
assign w1446 = ~w1443 & ~w1445;
assign w1447 = ~w1437 & w1441;
assign w1448 = w1437 & ~w1441;
assign w1449 = ~w1447 & ~w1448;
assign w1450 = w1442 & ~w1444;
assign w1451 = ~w1426 & ~w1431;
assign w1452 = ~w1450 & ~w1451;
assign w1453 = ~w1449 & ~w1452;
assign w1454 = ~w1446 & ~w1453;
assign w1455 = ~w1446 & ~w1452;
assign w1456 = A_844 & A_845;
assign w1457 = A_844 & ~A_845;
assign w1458 = ~A_844 & A_845;
assign w1459 = ~w1457 & ~w1458;
assign w1460 = (~w1456 & w1459) | (~w1456 & w13245) | (w1459 & w13245);
assign w1461 = A_841 & A_842;
assign w1462 = A_841 & ~A_842;
assign w1463 = ~A_841 & A_842;
assign w1464 = ~w1462 & ~w1463;
assign w1465 = (~w1461 & w1464) | (~w1461 & w13246) | (w1464 & w13246);
assign w1466 = ~w1460 & w1465;
assign w1467 = w1460 & ~w1465;
assign w1468 = ~w1466 & ~w1467;
assign w1469 = A_843 & ~w1462;
assign w1470 = ~w1463 & w1469;
assign w1471 = ~A_843 & ~w1464;
assign w1472 = ~w1470 & ~w1471;
assign w1473 = A_846 & ~w1457;
assign w1474 = ~w1458 & w1473;
assign w1475 = ~A_846 & ~w1459;
assign w1476 = ~w1474 & ~w1475;
assign w1477 = ~w1472 & ~w1476;
assign w1478 = ~w1468 & w1477;
assign w1479 = ~w1460 & ~w1465;
assign w1480 = ~w1478 & ~w1479;
assign w1481 = w1477 & w1468;
assign w1482 = ~w1468 & ~w1477;
assign w1483 = ~w1481 & ~w1482;
assign w1484 = ~w1480 & ~w1483;
assign w1485 = ~w1472 & w1476;
assign w1486 = w1472 & ~w1476;
assign w1487 = ~w1485 & ~w1486;
assign w1488 = ~w1449 & ~w1487;
assign w1489 = ~w1484 & w1488;
assign w1490 = ~w1455 & w1489;
assign w1491 = ~w1480 & ~w1487;
assign w1492 = ~w1483 & ~w1491;
assign w1493 = ~w1490 & ~w1492;
assign w1494 = ~w1483 & w1488;
assign w1495 = ~w1484 & w1494;
assign w1496 = ~w1455 & ~w1491;
assign w1497 = w1495 & w1496;
assign w1498 = (w1454 & w1493) | (w1454 & w13491) | (w1493 & w13491);
assign w1499 = ~w1490 & w1492;
assign w1500 = w1490 & ~w1492;
assign w1501 = ~w1499 & ~w1500;
assign w1502 = ~w1454 & ~w1501;
assign w1503 = ~w1484 & ~w1487;
assign w1504 = ~w1449 & ~w1455;
assign w1505 = ~w1503 & w1504;
assign w1506 = w1503 & ~w1504;
assign w1507 = ~w1505 & ~w1506;
assign w1508 = ~w1402 & ~w1405;
assign w1509 = ~w1367 & ~w1373;
assign w1510 = ~w1508 & w1509;
assign w1511 = w1508 & ~w1509;
assign w1512 = ~w1510 & ~w1511;
assign w1513 = ~w1507 & ~w1512;
assign w1514 = ~w1502 & w13492;
assign w1515 = (w1513 & w1502) | (w1513 & w13493) | (w1502 & w13493);
assign w1516 = ~w1514 & ~w1515;
assign w1517 = ~w1421 & ~w1516;
assign w1518 = ~w1502 & w13494;
assign w1519 = (~w1513 & w1502) | (~w1513 & w13683) | (w1502 & w13683);
assign w1520 = (w1421 & w1519) | (w1421 & w13495) | (w1519 & w13495);
assign w1521 = ~w1507 & w1512;
assign w1522 = w1507 & ~w1512;
assign w1523 = ~w1521 & ~w1522;
assign w1524 = ~w1243 & w1312;
assign w1525 = w1243 & ~w1312;
assign w1526 = ~w1524 & ~w1525;
assign w1527 = ~w1523 & ~w1526;
assign w1528 = ~w1527 & ~w1520;
assign w1529 = ~w1517 & w1528;
assign w1530 = ~w1517 & ~w1520;
assign w1531 = w1527 & ~w1530;
assign w1532 = (~w1339 & w1531) | (~w1339 & w13684) | (w1531 & w13684);
assign w1533 = w1527 & ~w1520;
assign w1534 = ~w1517 & w1533;
assign w1535 = ~w1527 & ~w1530;
assign w1536 = ~w1534 & ~w1535;
assign w1537 = (w1339 & w1535) | (w1339 & w13810) | (w1535 & w13810);
assign w1538 = ~w1523 & w1526;
assign w1539 = w1523 & ~w1526;
assign w1540 = ~w1538 & ~w1539;
assign w1541 = ~w961 & w1102;
assign w1542 = w961 & ~w1102;
assign w1543 = ~w1541 & ~w1542;
assign w1544 = ~w1540 & ~w1543;
assign w1545 = (~w1544 & w1536) | (~w1544 & w13685) | (w1536 & w13685);
assign w1546 = ~w1532 & w1545;
assign w1547 = (w1544 & w1537) | (w1544 & w13686) | (w1537 & w13686);
assign w1548 = ~w1546 & ~w1547;
assign w1549 = ~w1157 & ~w1548;
assign w1550 = (w1544 & w1536) | (w1544 & w13687) | (w1536 & w13687);
assign w1551 = ~w1532 & w1550;
assign w1552 = (~w1544 & w1537) | (~w1544 & w13688) | (w1537 & w13688);
assign w1553 = ~w1551 & ~w1552;
assign w1554 = w1157 & ~w1553;
assign w1555 = ~w1540 & w1543;
assign w1556 = w1540 & ~w1543;
assign w1557 = ~w1555 & ~w1556;
assign w1558 = ~w381 & w666;
assign w1559 = w381 & ~w666;
assign w1560 = ~w1558 & ~w1559;
assign w1561 = ~w1557 & ~w1560;
assign w1562 = (~w1561 & w1553) | (~w1561 & w13811) | (w1553 & w13811);
assign w1563 = ~w1549 & w1562;
assign w1564 = ~w1549 & ~w1554;
assign w1565 = w1561 & ~w1564;
assign w1566 = (~w777 & w1565) | (~w777 & w13812) | (w1565 & w13812);
assign w1567 = (w1561 & w1553) | (w1561 & w14055) | (w1553 & w14055);
assign w1568 = ~w1549 & w1567;
assign w1569 = ~w1561 & ~w1564;
assign w1570 = ~w1568 & ~w1569;
assign w1571 = (w777 & w1569) | (w777 & w14056) | (w1569 & w14056);
assign w1572 = ~A_469 & A_470;
assign w1573 = A_469 & ~A_470;
assign w1574 = A_471 & ~w1573;
assign w1575 = ~w1572 & w1574;
assign w1576 = ~w1572 & ~w1573;
assign w1577 = ~A_471 & ~w1576;
assign w1578 = ~w1575 & ~w1577;
assign w1579 = ~A_472 & A_473;
assign w1580 = A_472 & ~A_473;
assign w1581 = A_474 & ~w1580;
assign w1582 = ~w1579 & w1581;
assign w1583 = ~w1579 & ~w1580;
assign w1584 = ~A_474 & ~w1583;
assign w1585 = ~w1582 & ~w1584;
assign w1586 = ~w1578 & w1585;
assign w1587 = w1578 & ~w1585;
assign w1588 = ~w1586 & ~w1587;
assign w1589 = A_472 & A_473;
assign w1590 = (~w1589 & w1583) | (~w1589 & w13247) | (w1583 & w13247);
assign w1591 = A_469 & A_470;
assign w1592 = (~w1591 & w1576) | (~w1591 & w13248) | (w1576 & w13248);
assign w1593 = ~w1590 & w1592;
assign w1594 = w1590 & ~w1592;
assign w1595 = ~w1593 & ~w1594;
assign w1596 = ~w1578 & ~w1585;
assign w1597 = ~w1595 & w1596;
assign w1598 = ~w1590 & ~w1592;
assign w1599 = ~w1597 & ~w1598;
assign w1600 = w1596 & w1595;
assign w1601 = ~w1595 & ~w1596;
assign w1602 = ~w1600 & ~w1601;
assign w1603 = ~w1599 & ~w1602;
assign w1604 = ~w1588 & ~w1603;
assign w1605 = ~A_466 & A_467;
assign w1606 = A_466 & ~A_467;
assign w1607 = A_468 & ~w1606;
assign w1608 = ~w1605 & w1607;
assign w1609 = ~w1605 & ~w1606;
assign w1610 = ~A_468 & ~w1609;
assign w1611 = ~w1608 & ~w1610;
assign w1612 = ~A_463 & A_464;
assign w1613 = A_463 & ~A_464;
assign w1614 = A_465 & ~w1613;
assign w1615 = ~w1612 & w1614;
assign w1616 = ~w1612 & ~w1613;
assign w1617 = ~A_465 & ~w1616;
assign w1618 = ~w1615 & ~w1617;
assign w1619 = ~w1611 & w1618;
assign w1620 = w1611 & ~w1618;
assign w1621 = ~w1619 & ~w1620;
assign w1622 = A_466 & A_467;
assign w1623 = (~w1622 & w1609) | (~w1622 & w13249) | (w1609 & w13249);
assign w1624 = A_463 & A_464;
assign w1625 = (~w1624 & w1616) | (~w1624 & w13250) | (w1616 & w13250);
assign w1626 = w1623 & ~w1625;
assign w1627 = ~w1623 & w1625;
assign w1628 = ~w1611 & ~w1618;
assign w1629 = w1628 & w1630;
assign w1630 = ~w1626 & ~w1627;
assign w1631 = ~w1628 & ~w1630;
assign w1632 = ~w1629 & ~w1631;
assign w1633 = w1628 & ~w1630;
assign w1634 = ~w1623 & ~w1625;
assign w1635 = ~w1633 & ~w1634;
assign w1636 = ~w1632 & ~w1635;
assign w1637 = ~w1621 & ~w1636;
assign w1638 = ~w1604 & w1637;
assign w1639 = w1604 & ~w1637;
assign w1640 = ~w1638 & ~w1639;
assign w1641 = ~A_481 & A_482;
assign w1642 = A_481 & ~A_482;
assign w1643 = A_483 & ~w1642;
assign w1644 = ~w1641 & w1643;
assign w1645 = ~w1641 & ~w1642;
assign w1646 = ~A_483 & ~w1645;
assign w1647 = ~w1644 & ~w1646;
assign w1648 = ~A_484 & A_485;
assign w1649 = A_484 & ~A_485;
assign w1650 = A_486 & ~w1649;
assign w1651 = ~w1648 & w1650;
assign w1652 = ~w1648 & ~w1649;
assign w1653 = ~A_486 & ~w1652;
assign w1654 = ~w1651 & ~w1653;
assign w1655 = ~w1647 & w1654;
assign w1656 = w1647 & ~w1654;
assign w1657 = ~w1655 & ~w1656;
assign w1658 = A_484 & A_485;
assign w1659 = (~w1658 & w1652) | (~w1658 & w13251) | (w1652 & w13251);
assign w1660 = A_481 & A_482;
assign w1661 = (~w1660 & w1645) | (~w1660 & w13252) | (w1645 & w13252);
assign w1662 = ~w1659 & w1661;
assign w1663 = w1659 & ~w1661;
assign w1664 = ~w1662 & ~w1663;
assign w1665 = ~w1647 & ~w1654;
assign w1666 = ~w1664 & w1665;
assign w1667 = ~w1659 & ~w1661;
assign w1668 = ~w1666 & ~w1667;
assign w1669 = w1665 & w1664;
assign w1670 = ~w1664 & ~w1665;
assign w1671 = ~w1669 & ~w1670;
assign w1672 = ~w1668 & ~w1671;
assign w1673 = ~w1657 & ~w1672;
assign w1674 = ~A_475 & A_476;
assign w1675 = A_475 & ~A_476;
assign w1676 = A_477 & ~w1675;
assign w1677 = ~w1674 & w1676;
assign w1678 = ~w1674 & ~w1675;
assign w1679 = ~A_477 & ~w1678;
assign w1680 = ~w1677 & ~w1679;
assign w1681 = ~A_478 & A_479;
assign w1682 = A_478 & ~A_479;
assign w1683 = A_480 & ~w1682;
assign w1684 = ~w1681 & w1683;
assign w1685 = ~w1681 & ~w1682;
assign w1686 = ~A_480 & ~w1685;
assign w1687 = ~w1684 & ~w1686;
assign w1688 = ~w1680 & w1687;
assign w1689 = w1680 & ~w1687;
assign w1690 = ~w1688 & ~w1689;
assign w1691 = A_478 & A_479;
assign w1692 = (~w1691 & w1685) | (~w1691 & w13253) | (w1685 & w13253);
assign w1693 = A_475 & A_476;
assign w1694 = (~w1693 & w1678) | (~w1693 & w13254) | (w1678 & w13254);
assign w1695 = ~w1692 & w1694;
assign w1696 = w1692 & ~w1694;
assign w1697 = ~w1695 & ~w1696;
assign w1698 = ~w1680 & ~w1687;
assign w1699 = ~w1697 & w1698;
assign w1700 = ~w1692 & ~w1694;
assign w1701 = ~w1699 & ~w1700;
assign w1702 = w1698 & w1697;
assign w1703 = ~w1697 & ~w1698;
assign w1704 = ~w1702 & ~w1703;
assign w1705 = ~w1701 & ~w1704;
assign w1706 = ~w1690 & ~w1705;
assign w1707 = ~w1673 & w1706;
assign w1708 = w1673 & ~w1706;
assign w1709 = ~w1707 & ~w1708;
assign w1710 = ~w1640 & w1709;
assign w1711 = w1640 & ~w1709;
assign w1712 = ~w1710 & ~w1711;
assign w1713 = ~A_505 & A_506;
assign w1714 = A_505 & ~A_506;
assign w1715 = A_507 & ~w1714;
assign w1716 = ~w1713 & w1715;
assign w1717 = ~w1713 & ~w1714;
assign w1718 = ~A_507 & ~w1717;
assign w1719 = ~w1716 & ~w1718;
assign w1720 = ~A_508 & A_509;
assign w1721 = A_508 & ~A_509;
assign w1722 = A_510 & ~w1721;
assign w1723 = ~w1720 & w1722;
assign w1724 = ~w1720 & ~w1721;
assign w1725 = ~A_510 & ~w1724;
assign w1726 = ~w1723 & ~w1725;
assign w1727 = ~w1719 & w1726;
assign w1728 = w1719 & ~w1726;
assign w1729 = ~w1727 & ~w1728;
assign w1730 = A_508 & A_509;
assign w1731 = (~w1730 & w1724) | (~w1730 & w13255) | (w1724 & w13255);
assign w1732 = A_505 & A_506;
assign w1733 = (~w1732 & w1717) | (~w1732 & w13256) | (w1717 & w13256);
assign w1734 = ~w1731 & w1733;
assign w1735 = w1731 & ~w1733;
assign w1736 = ~w1734 & ~w1735;
assign w1737 = ~w1719 & ~w1726;
assign w1738 = ~w1736 & w1737;
assign w1739 = ~w1731 & ~w1733;
assign w1740 = ~w1738 & ~w1739;
assign w1741 = w1737 & w1736;
assign w1742 = ~w1736 & ~w1737;
assign w1743 = ~w1741 & ~w1742;
assign w1744 = ~w1740 & ~w1743;
assign w1745 = ~w1729 & ~w1744;
assign w1746 = ~A_499 & A_500;
assign w1747 = A_499 & ~A_500;
assign w1748 = A_501 & ~w1747;
assign w1749 = ~w1746 & w1748;
assign w1750 = ~w1746 & ~w1747;
assign w1751 = ~A_501 & ~w1750;
assign w1752 = ~w1749 & ~w1751;
assign w1753 = ~A_502 & A_503;
assign w1754 = A_502 & ~A_503;
assign w1755 = A_504 & ~w1754;
assign w1756 = ~w1753 & w1755;
assign w1757 = ~w1753 & ~w1754;
assign w1758 = ~A_504 & ~w1757;
assign w1759 = ~w1756 & ~w1758;
assign w1760 = ~w1752 & w1759;
assign w1761 = w1752 & ~w1759;
assign w1762 = ~w1760 & ~w1761;
assign w1763 = A_502 & A_503;
assign w1764 = (~w1763 & w1757) | (~w1763 & w13257) | (w1757 & w13257);
assign w1765 = A_499 & A_500;
assign w1766 = (~w1765 & w1750) | (~w1765 & w13258) | (w1750 & w13258);
assign w1767 = ~w1764 & w1766;
assign w1768 = w1764 & ~w1766;
assign w1769 = ~w1767 & ~w1768;
assign w1770 = ~w1752 & ~w1759;
assign w1771 = ~w1769 & w1770;
assign w1772 = ~w1764 & ~w1766;
assign w1773 = ~w1771 & ~w1772;
assign w1774 = w1770 & w1769;
assign w1775 = ~w1769 & ~w1770;
assign w1776 = ~w1774 & ~w1775;
assign w1777 = ~w1773 & ~w1776;
assign w1778 = ~w1762 & ~w1777;
assign w1779 = ~w1745 & w1778;
assign w1780 = w1745 & ~w1778;
assign w1781 = ~w1779 & ~w1780;
assign w1782 = ~A_493 & A_494;
assign w1783 = A_493 & ~A_494;
assign w1784 = A_495 & ~w1783;
assign w1785 = ~w1782 & w1784;
assign w1786 = ~w1782 & ~w1783;
assign w1787 = ~A_495 & ~w1786;
assign w1788 = ~w1785 & ~w1787;
assign w1789 = ~A_496 & A_497;
assign w1790 = A_496 & ~A_497;
assign w1791 = A_498 & ~w1790;
assign w1792 = ~w1789 & w1791;
assign w1793 = ~w1789 & ~w1790;
assign w1794 = ~A_498 & ~w1793;
assign w1795 = ~w1792 & ~w1794;
assign w1796 = ~w1788 & w1795;
assign w1797 = w1788 & ~w1795;
assign w1798 = ~w1796 & ~w1797;
assign w1799 = A_496 & A_497;
assign w1800 = (~w1799 & w1793) | (~w1799 & w13259) | (w1793 & w13259);
assign w1801 = A_493 & A_494;
assign w1802 = (~w1801 & w1786) | (~w1801 & w13260) | (w1786 & w13260);
assign w1803 = ~w1800 & w1802;
assign w1804 = w1800 & ~w1802;
assign w1805 = ~w1803 & ~w1804;
assign w1806 = ~w1788 & ~w1795;
assign w1807 = ~w1805 & w1806;
assign w1808 = ~w1800 & ~w1802;
assign w1809 = ~w1807 & ~w1808;
assign w1810 = w1806 & w1805;
assign w1811 = ~w1805 & ~w1806;
assign w1812 = ~w1810 & ~w1811;
assign w1813 = ~w1809 & ~w1812;
assign w1814 = ~w1798 & ~w1813;
assign w1815 = ~A_487 & A_488;
assign w1816 = A_487 & ~A_488;
assign w1817 = A_489 & ~w1816;
assign w1818 = ~w1815 & w1817;
assign w1819 = ~w1815 & ~w1816;
assign w1820 = ~A_489 & ~w1819;
assign w1821 = ~w1818 & ~w1820;
assign w1822 = ~A_490 & A_491;
assign w1823 = A_490 & ~A_491;
assign w1824 = A_492 & ~w1823;
assign w1825 = ~w1822 & w1824;
assign w1826 = ~w1822 & ~w1823;
assign w1827 = ~A_492 & ~w1826;
assign w1828 = ~w1825 & ~w1827;
assign w1829 = ~w1821 & w1828;
assign w1830 = w1821 & ~w1828;
assign w1831 = ~w1829 & ~w1830;
assign w1832 = A_490 & A_491;
assign w1833 = (~w1832 & w1826) | (~w1832 & w13261) | (w1826 & w13261);
assign w1834 = A_487 & A_488;
assign w1835 = (~w1834 & w1819) | (~w1834 & w13262) | (w1819 & w13262);
assign w1836 = ~w1833 & w1835;
assign w1837 = w1833 & ~w1835;
assign w1838 = ~w1836 & ~w1837;
assign w1839 = ~w1821 & ~w1828;
assign w1840 = ~w1838 & w1839;
assign w1841 = ~w1833 & ~w1835;
assign w1842 = ~w1840 & ~w1841;
assign w1843 = w1839 & w1838;
assign w1844 = ~w1838 & ~w1839;
assign w1845 = ~w1843 & ~w1844;
assign w1846 = ~w1842 & ~w1845;
assign w1847 = ~w1831 & ~w1846;
assign w1848 = ~w1814 & w1847;
assign w1849 = w1814 & ~w1847;
assign w1850 = ~w1848 & ~w1849;
assign w1851 = ~w1781 & w1850;
assign w1852 = w1781 & ~w1850;
assign w1853 = ~w1851 & ~w1852;
assign w1854 = ~w1712 & w1853;
assign w1855 = w1712 & ~w1853;
assign w1856 = ~w1854 & ~w1855;
assign w1857 = ~A_553 & A_554;
assign w1858 = A_553 & ~A_554;
assign w1859 = A_555 & ~w1858;
assign w1860 = ~w1857 & w1859;
assign w1861 = ~w1857 & ~w1858;
assign w1862 = ~A_555 & ~w1861;
assign w1863 = ~w1860 & ~w1862;
assign w1864 = ~A_556 & A_557;
assign w1865 = A_556 & ~A_557;
assign w1866 = A_558 & ~w1865;
assign w1867 = ~w1864 & w1866;
assign w1868 = ~w1864 & ~w1865;
assign w1869 = ~A_558 & ~w1868;
assign w1870 = ~w1867 & ~w1869;
assign w1871 = ~w1863 & w1870;
assign w1872 = w1863 & ~w1870;
assign w1873 = ~w1871 & ~w1872;
assign w1874 = A_556 & A_557;
assign w1875 = (~w1874 & w1868) | (~w1874 & w13263) | (w1868 & w13263);
assign w1876 = A_553 & A_554;
assign w1877 = (~w1876 & w1861) | (~w1876 & w13264) | (w1861 & w13264);
assign w1878 = ~w1875 & w1877;
assign w1879 = w1875 & ~w1877;
assign w1880 = ~w1878 & ~w1879;
assign w1881 = ~w1863 & ~w1870;
assign w1882 = ~w1880 & w1881;
assign w1883 = ~w1875 & ~w1877;
assign w1884 = ~w1882 & ~w1883;
assign w1885 = w1881 & w1880;
assign w1886 = ~w1880 & ~w1881;
assign w1887 = ~w1885 & ~w1886;
assign w1888 = ~w1884 & ~w1887;
assign w1889 = ~w1873 & ~w1888;
assign w1890 = ~A_547 & A_548;
assign w1891 = A_547 & ~A_548;
assign w1892 = A_549 & ~w1891;
assign w1893 = ~w1890 & w1892;
assign w1894 = ~w1890 & ~w1891;
assign w1895 = ~A_549 & ~w1894;
assign w1896 = ~w1893 & ~w1895;
assign w1897 = ~A_550 & A_551;
assign w1898 = A_550 & ~A_551;
assign w1899 = A_552 & ~w1898;
assign w1900 = ~w1897 & w1899;
assign w1901 = ~w1897 & ~w1898;
assign w1902 = ~A_552 & ~w1901;
assign w1903 = ~w1900 & ~w1902;
assign w1904 = ~w1896 & w1903;
assign w1905 = w1896 & ~w1903;
assign w1906 = ~w1904 & ~w1905;
assign w1907 = A_550 & A_551;
assign w1908 = (~w1907 & w1901) | (~w1907 & w13265) | (w1901 & w13265);
assign w1909 = A_547 & A_548;
assign w1910 = (~w1909 & w1894) | (~w1909 & w13266) | (w1894 & w13266);
assign w1911 = ~w1908 & w1910;
assign w1912 = w1908 & ~w1910;
assign w1913 = ~w1911 & ~w1912;
assign w1914 = ~w1896 & ~w1903;
assign w1915 = ~w1913 & w1914;
assign w1916 = ~w1908 & ~w1910;
assign w1917 = ~w1915 & ~w1916;
assign w1918 = w1914 & w1913;
assign w1919 = ~w1913 & ~w1914;
assign w1920 = ~w1918 & ~w1919;
assign w1921 = ~w1917 & ~w1920;
assign w1922 = ~w1906 & ~w1921;
assign w1923 = ~w1889 & w1922;
assign w1924 = w1889 & ~w1922;
assign w1925 = ~w1923 & ~w1924;
assign w1926 = ~A_541 & A_542;
assign w1927 = A_541 & ~A_542;
assign w1928 = A_543 & ~w1927;
assign w1929 = ~w1926 & w1928;
assign w1930 = ~w1926 & ~w1927;
assign w1931 = ~A_543 & ~w1930;
assign w1932 = ~w1929 & ~w1931;
assign w1933 = ~A_544 & A_545;
assign w1934 = A_544 & ~A_545;
assign w1935 = A_546 & ~w1934;
assign w1936 = ~w1933 & w1935;
assign w1937 = ~w1933 & ~w1934;
assign w1938 = ~A_546 & ~w1937;
assign w1939 = ~w1936 & ~w1938;
assign w1940 = ~w1932 & w1939;
assign w1941 = w1932 & ~w1939;
assign w1942 = ~w1940 & ~w1941;
assign w1943 = A_544 & A_545;
assign w1944 = (~w1943 & w1937) | (~w1943 & w13267) | (w1937 & w13267);
assign w1945 = A_541 & A_542;
assign w1946 = (~w1945 & w1930) | (~w1945 & w13268) | (w1930 & w13268);
assign w1947 = ~w1944 & w1946;
assign w1948 = w1944 & ~w1946;
assign w1949 = ~w1947 & ~w1948;
assign w1950 = ~w1932 & ~w1939;
assign w1951 = ~w1949 & w1950;
assign w1952 = ~w1944 & ~w1946;
assign w1953 = ~w1951 & ~w1952;
assign w1954 = w1950 & w1949;
assign w1955 = ~w1949 & ~w1950;
assign w1956 = ~w1954 & ~w1955;
assign w1957 = ~w1953 & ~w1956;
assign w1958 = ~w1942 & ~w1957;
assign w1959 = ~A_535 & A_536;
assign w1960 = A_535 & ~A_536;
assign w1961 = A_537 & ~w1960;
assign w1962 = ~w1959 & w1961;
assign w1963 = ~w1959 & ~w1960;
assign w1964 = ~A_537 & ~w1963;
assign w1965 = ~w1962 & ~w1964;
assign w1966 = ~A_538 & A_539;
assign w1967 = A_538 & ~A_539;
assign w1968 = A_540 & ~w1967;
assign w1969 = ~w1966 & w1968;
assign w1970 = ~w1966 & ~w1967;
assign w1971 = ~A_540 & ~w1970;
assign w1972 = ~w1969 & ~w1971;
assign w1973 = ~w1965 & w1972;
assign w1974 = w1965 & ~w1972;
assign w1975 = ~w1973 & ~w1974;
assign w1976 = A_538 & A_539;
assign w1977 = (~w1976 & w1970) | (~w1976 & w13269) | (w1970 & w13269);
assign w1978 = A_535 & A_536;
assign w1979 = (~w1978 & w1963) | (~w1978 & w13270) | (w1963 & w13270);
assign w1980 = ~w1977 & w1979;
assign w1981 = w1977 & ~w1979;
assign w1982 = ~w1980 & ~w1981;
assign w1983 = ~w1965 & ~w1972;
assign w1984 = ~w1982 & w1983;
assign w1985 = ~w1977 & ~w1979;
assign w1986 = ~w1984 & ~w1985;
assign w1987 = w1983 & w1982;
assign w1988 = ~w1982 & ~w1983;
assign w1989 = ~w1987 & ~w1988;
assign w1990 = ~w1986 & ~w1989;
assign w1991 = ~w1975 & ~w1990;
assign w1992 = ~w1958 & w1991;
assign w1993 = w1958 & ~w1991;
assign w1994 = ~w1992 & ~w1993;
assign w1995 = ~w1925 & w1994;
assign w1996 = w1925 & ~w1994;
assign w1997 = ~w1995 & ~w1996;
assign w1998 = ~A_529 & A_530;
assign w1999 = A_529 & ~A_530;
assign w2000 = A_531 & ~w1999;
assign w2001 = ~w1998 & w2000;
assign w2002 = ~w1998 & ~w1999;
assign w2003 = ~A_531 & ~w2002;
assign w2004 = ~w2001 & ~w2003;
assign w2005 = ~A_532 & A_533;
assign w2006 = A_532 & ~A_533;
assign w2007 = A_534 & ~w2006;
assign w2008 = ~w2005 & w2007;
assign w2009 = ~w2005 & ~w2006;
assign w2010 = ~A_534 & ~w2009;
assign w2011 = ~w2008 & ~w2010;
assign w2012 = ~w2004 & w2011;
assign w2013 = w2004 & ~w2011;
assign w2014 = ~w2012 & ~w2013;
assign w2015 = A_532 & A_533;
assign w2016 = (~w2015 & w2009) | (~w2015 & w13271) | (w2009 & w13271);
assign w2017 = A_529 & A_530;
assign w2018 = (~w2017 & w2002) | (~w2017 & w13272) | (w2002 & w13272);
assign w2019 = ~w2016 & w2018;
assign w2020 = w2016 & ~w2018;
assign w2021 = ~w2019 & ~w2020;
assign w2022 = ~w2004 & ~w2011;
assign w2023 = ~w2021 & w2022;
assign w2024 = ~w2016 & ~w2018;
assign w2025 = ~w2023 & ~w2024;
assign w2026 = w2022 & w2021;
assign w2027 = ~w2021 & ~w2022;
assign w2028 = ~w2026 & ~w2027;
assign w2029 = ~w2025 & ~w2028;
assign w2030 = ~w2014 & ~w2029;
assign w2031 = ~A_523 & A_524;
assign w2032 = A_523 & ~A_524;
assign w2033 = A_525 & ~w2032;
assign w2034 = ~w2031 & w2033;
assign w2035 = ~w2031 & ~w2032;
assign w2036 = ~A_525 & ~w2035;
assign w2037 = ~w2034 & ~w2036;
assign w2038 = ~A_526 & A_527;
assign w2039 = A_526 & ~A_527;
assign w2040 = A_528 & ~w2039;
assign w2041 = ~w2038 & w2040;
assign w2042 = ~w2038 & ~w2039;
assign w2043 = ~A_528 & ~w2042;
assign w2044 = ~w2041 & ~w2043;
assign w2045 = ~w2037 & w2044;
assign w2046 = w2037 & ~w2044;
assign w2047 = ~w2045 & ~w2046;
assign w2048 = A_526 & A_527;
assign w2049 = (~w2048 & w2042) | (~w2048 & w13273) | (w2042 & w13273);
assign w2050 = A_523 & A_524;
assign w2051 = (~w2050 & w2035) | (~w2050 & w13274) | (w2035 & w13274);
assign w2052 = ~w2049 & w2051;
assign w2053 = w2049 & ~w2051;
assign w2054 = ~w2052 & ~w2053;
assign w2055 = ~w2037 & ~w2044;
assign w2056 = ~w2054 & w2055;
assign w2057 = ~w2049 & ~w2051;
assign w2058 = ~w2056 & ~w2057;
assign w2059 = w2055 & w2054;
assign w2060 = ~w2054 & ~w2055;
assign w2061 = ~w2059 & ~w2060;
assign w2062 = ~w2058 & ~w2061;
assign w2063 = ~w2047 & ~w2062;
assign w2064 = ~w2030 & w2063;
assign w2065 = w2030 & ~w2063;
assign w2066 = ~w2064 & ~w2065;
assign w2067 = ~A_517 & A_518;
assign w2068 = A_517 & ~A_518;
assign w2069 = A_519 & ~w2068;
assign w2070 = ~w2067 & w2069;
assign w2071 = ~w2067 & ~w2068;
assign w2072 = ~A_519 & ~w2071;
assign w2073 = ~w2070 & ~w2072;
assign w2074 = ~A_520 & A_521;
assign w2075 = A_520 & ~A_521;
assign w2076 = A_522 & ~w2075;
assign w2077 = ~w2074 & w2076;
assign w2078 = ~w2074 & ~w2075;
assign w2079 = ~A_522 & ~w2078;
assign w2080 = ~w2077 & ~w2079;
assign w2081 = ~w2073 & w2080;
assign w2082 = w2073 & ~w2080;
assign w2083 = ~w2081 & ~w2082;
assign w2084 = A_520 & A_521;
assign w2085 = (~w2084 & w2078) | (~w2084 & w13275) | (w2078 & w13275);
assign w2086 = A_517 & A_518;
assign w2087 = (~w2086 & w2071) | (~w2086 & w13276) | (w2071 & w13276);
assign w2088 = ~w2085 & w2087;
assign w2089 = w2085 & ~w2087;
assign w2090 = ~w2088 & ~w2089;
assign w2091 = ~w2073 & ~w2080;
assign w2092 = ~w2090 & w2091;
assign w2093 = ~w2085 & ~w2087;
assign w2094 = ~w2092 & ~w2093;
assign w2095 = w2091 & w2090;
assign w2096 = ~w2090 & ~w2091;
assign w2097 = ~w2095 & ~w2096;
assign w2098 = ~w2094 & ~w2097;
assign w2099 = ~w2083 & ~w2098;
assign w2100 = ~A_511 & A_512;
assign w2101 = A_511 & ~A_512;
assign w2102 = A_513 & ~w2101;
assign w2103 = ~w2100 & w2102;
assign w2104 = ~w2100 & ~w2101;
assign w2105 = ~A_513 & ~w2104;
assign w2106 = ~w2103 & ~w2105;
assign w2107 = ~A_514 & A_515;
assign w2108 = A_514 & ~A_515;
assign w2109 = A_516 & ~w2108;
assign w2110 = ~w2107 & w2109;
assign w2111 = ~w2107 & ~w2108;
assign w2112 = ~A_516 & ~w2111;
assign w2113 = ~w2110 & ~w2112;
assign w2114 = ~w2106 & w2113;
assign w2115 = w2106 & ~w2113;
assign w2116 = ~w2114 & ~w2115;
assign w2117 = A_514 & A_515;
assign w2118 = (~w2117 & w2111) | (~w2117 & w13277) | (w2111 & w13277);
assign w2119 = A_511 & A_512;
assign w2120 = (~w2119 & w2104) | (~w2119 & w13278) | (w2104 & w13278);
assign w2121 = ~w2118 & w2120;
assign w2122 = w2118 & ~w2120;
assign w2123 = ~w2121 & ~w2122;
assign w2124 = ~w2106 & ~w2113;
assign w2125 = ~w2123 & w2124;
assign w2126 = ~w2118 & ~w2120;
assign w2127 = ~w2125 & ~w2126;
assign w2128 = w2124 & w2123;
assign w2129 = ~w2123 & ~w2124;
assign w2130 = ~w2128 & ~w2129;
assign w2131 = ~w2127 & ~w2130;
assign w2132 = ~w2116 & ~w2131;
assign w2133 = ~w2099 & w2132;
assign w2134 = w2099 & ~w2132;
assign w2135 = ~w2133 & ~w2134;
assign w2136 = ~w2066 & w2135;
assign w2137 = w2066 & ~w2135;
assign w2138 = ~w2136 & ~w2137;
assign w2139 = ~w1997 & w2138;
assign w2140 = w1997 & ~w2138;
assign w2141 = ~w2139 & ~w2140;
assign w2142 = ~w1856 & w2141;
assign w2143 = w1856 & ~w2141;
assign w2144 = ~w2142 & ~w2143;
assign w2145 = ~A_649 & A_650;
assign w2146 = A_649 & ~A_650;
assign w2147 = A_651 & ~w2146;
assign w2148 = ~w2145 & w2147;
assign w2149 = ~w2145 & ~w2146;
assign w2150 = ~A_651 & ~w2149;
assign w2151 = ~w2148 & ~w2150;
assign w2152 = ~A_652 & A_653;
assign w2153 = A_652 & ~A_653;
assign w2154 = A_654 & ~w2153;
assign w2155 = ~w2152 & w2154;
assign w2156 = ~w2152 & ~w2153;
assign w2157 = ~A_654 & ~w2156;
assign w2158 = ~w2155 & ~w2157;
assign w2159 = ~w2151 & w2158;
assign w2160 = w2151 & ~w2158;
assign w2161 = ~w2159 & ~w2160;
assign w2162 = A_652 & A_653;
assign w2163 = (~w2162 & w2156) | (~w2162 & w13279) | (w2156 & w13279);
assign w2164 = A_649 & A_650;
assign w2165 = (~w2164 & w2149) | (~w2164 & w13280) | (w2149 & w13280);
assign w2166 = ~w2163 & w2165;
assign w2167 = w2163 & ~w2165;
assign w2168 = ~w2166 & ~w2167;
assign w2169 = ~w2151 & ~w2158;
assign w2170 = ~w2168 & w2169;
assign w2171 = ~w2163 & ~w2165;
assign w2172 = ~w2170 & ~w2171;
assign w2173 = w2169 & w2168;
assign w2174 = ~w2168 & ~w2169;
assign w2175 = ~w2173 & ~w2174;
assign w2176 = ~w2172 & ~w2175;
assign w2177 = ~w2161 & ~w2176;
assign w2178 = ~A_643 & A_644;
assign w2179 = A_643 & ~A_644;
assign w2180 = A_645 & ~w2179;
assign w2181 = ~w2178 & w2180;
assign w2182 = ~w2178 & ~w2179;
assign w2183 = ~A_645 & ~w2182;
assign w2184 = ~w2181 & ~w2183;
assign w2185 = ~A_646 & A_647;
assign w2186 = A_646 & ~A_647;
assign w2187 = A_648 & ~w2186;
assign w2188 = ~w2185 & w2187;
assign w2189 = ~w2185 & ~w2186;
assign w2190 = ~A_648 & ~w2189;
assign w2191 = ~w2188 & ~w2190;
assign w2192 = ~w2184 & w2191;
assign w2193 = w2184 & ~w2191;
assign w2194 = ~w2192 & ~w2193;
assign w2195 = A_646 & A_647;
assign w2196 = (~w2195 & w2189) | (~w2195 & w13281) | (w2189 & w13281);
assign w2197 = A_643 & A_644;
assign w2198 = (~w2197 & w2182) | (~w2197 & w13282) | (w2182 & w13282);
assign w2199 = ~w2196 & w2198;
assign w2200 = w2196 & ~w2198;
assign w2201 = ~w2199 & ~w2200;
assign w2202 = ~w2184 & ~w2191;
assign w2203 = ~w2201 & w2202;
assign w2204 = ~w2196 & ~w2198;
assign w2205 = ~w2203 & ~w2204;
assign w2206 = w2202 & w2201;
assign w2207 = ~w2201 & ~w2202;
assign w2208 = ~w2206 & ~w2207;
assign w2209 = ~w2205 & ~w2208;
assign w2210 = ~w2194 & ~w2209;
assign w2211 = ~w2177 & w2210;
assign w2212 = w2177 & ~w2210;
assign w2213 = ~w2211 & ~w2212;
assign w2214 = ~A_637 & A_638;
assign w2215 = A_637 & ~A_638;
assign w2216 = A_639 & ~w2215;
assign w2217 = ~w2214 & w2216;
assign w2218 = ~w2214 & ~w2215;
assign w2219 = ~A_639 & ~w2218;
assign w2220 = ~w2217 & ~w2219;
assign w2221 = ~A_640 & A_641;
assign w2222 = A_640 & ~A_641;
assign w2223 = A_642 & ~w2222;
assign w2224 = ~w2221 & w2223;
assign w2225 = ~w2221 & ~w2222;
assign w2226 = ~A_642 & ~w2225;
assign w2227 = ~w2224 & ~w2226;
assign w2228 = ~w2220 & w2227;
assign w2229 = w2220 & ~w2227;
assign w2230 = ~w2228 & ~w2229;
assign w2231 = A_640 & A_641;
assign w2232 = (~w2231 & w2225) | (~w2231 & w13283) | (w2225 & w13283);
assign w2233 = A_637 & A_638;
assign w2234 = (~w2233 & w2218) | (~w2233 & w13284) | (w2218 & w13284);
assign w2235 = ~w2232 & w2234;
assign w2236 = w2232 & ~w2234;
assign w2237 = ~w2235 & ~w2236;
assign w2238 = ~w2220 & ~w2227;
assign w2239 = ~w2237 & w2238;
assign w2240 = ~w2232 & ~w2234;
assign w2241 = ~w2239 & ~w2240;
assign w2242 = w2238 & w2237;
assign w2243 = ~w2237 & ~w2238;
assign w2244 = ~w2242 & ~w2243;
assign w2245 = ~w2241 & ~w2244;
assign w2246 = ~w2230 & ~w2245;
assign w2247 = ~A_631 & A_632;
assign w2248 = A_631 & ~A_632;
assign w2249 = A_633 & ~w2248;
assign w2250 = ~w2247 & w2249;
assign w2251 = ~w2247 & ~w2248;
assign w2252 = ~A_633 & ~w2251;
assign w2253 = ~w2250 & ~w2252;
assign w2254 = ~A_634 & A_635;
assign w2255 = A_634 & ~A_635;
assign w2256 = A_636 & ~w2255;
assign w2257 = ~w2254 & w2256;
assign w2258 = ~w2254 & ~w2255;
assign w2259 = ~A_636 & ~w2258;
assign w2260 = ~w2257 & ~w2259;
assign w2261 = ~w2253 & w2260;
assign w2262 = w2253 & ~w2260;
assign w2263 = ~w2261 & ~w2262;
assign w2264 = A_634 & A_635;
assign w2265 = (~w2264 & w2258) | (~w2264 & w13285) | (w2258 & w13285);
assign w2266 = A_631 & A_632;
assign w2267 = (~w2266 & w2251) | (~w2266 & w13286) | (w2251 & w13286);
assign w2268 = ~w2265 & w2267;
assign w2269 = w2265 & ~w2267;
assign w2270 = ~w2268 & ~w2269;
assign w2271 = ~w2253 & ~w2260;
assign w2272 = ~w2270 & w2271;
assign w2273 = ~w2265 & ~w2267;
assign w2274 = ~w2272 & ~w2273;
assign w2275 = w2271 & w2270;
assign w2276 = ~w2270 & ~w2271;
assign w2277 = ~w2275 & ~w2276;
assign w2278 = ~w2274 & ~w2277;
assign w2279 = ~w2263 & ~w2278;
assign w2280 = ~w2246 & w2279;
assign w2281 = w2246 & ~w2279;
assign w2282 = ~w2280 & ~w2281;
assign w2283 = ~w2213 & w2282;
assign w2284 = w2213 & ~w2282;
assign w2285 = ~w2283 & ~w2284;
assign w2286 = ~A_625 & A_626;
assign w2287 = A_625 & ~A_626;
assign w2288 = A_627 & ~w2287;
assign w2289 = ~w2286 & w2288;
assign w2290 = ~w2286 & ~w2287;
assign w2291 = ~A_627 & ~w2290;
assign w2292 = ~w2289 & ~w2291;
assign w2293 = ~A_628 & A_629;
assign w2294 = A_628 & ~A_629;
assign w2295 = A_630 & ~w2294;
assign w2296 = ~w2293 & w2295;
assign w2297 = ~w2293 & ~w2294;
assign w2298 = ~A_630 & ~w2297;
assign w2299 = ~w2296 & ~w2298;
assign w2300 = ~w2292 & w2299;
assign w2301 = w2292 & ~w2299;
assign w2302 = ~w2300 & ~w2301;
assign w2303 = A_628 & A_629;
assign w2304 = (~w2303 & w2297) | (~w2303 & w13287) | (w2297 & w13287);
assign w2305 = A_625 & A_626;
assign w2306 = (~w2305 & w2290) | (~w2305 & w13288) | (w2290 & w13288);
assign w2307 = ~w2304 & w2306;
assign w2308 = w2304 & ~w2306;
assign w2309 = ~w2307 & ~w2308;
assign w2310 = ~w2292 & ~w2299;
assign w2311 = ~w2309 & w2310;
assign w2312 = ~w2304 & ~w2306;
assign w2313 = ~w2311 & ~w2312;
assign w2314 = w2310 & w2309;
assign w2315 = ~w2309 & ~w2310;
assign w2316 = ~w2314 & ~w2315;
assign w2317 = ~w2313 & ~w2316;
assign w2318 = ~w2302 & ~w2317;
assign w2319 = ~A_619 & A_620;
assign w2320 = A_619 & ~A_620;
assign w2321 = A_621 & ~w2320;
assign w2322 = ~w2319 & w2321;
assign w2323 = ~w2319 & ~w2320;
assign w2324 = ~A_621 & ~w2323;
assign w2325 = ~w2322 & ~w2324;
assign w2326 = ~A_622 & A_623;
assign w2327 = A_622 & ~A_623;
assign w2328 = A_624 & ~w2327;
assign w2329 = ~w2326 & w2328;
assign w2330 = ~w2326 & ~w2327;
assign w2331 = ~A_624 & ~w2330;
assign w2332 = ~w2329 & ~w2331;
assign w2333 = ~w2325 & w2332;
assign w2334 = w2325 & ~w2332;
assign w2335 = ~w2333 & ~w2334;
assign w2336 = A_622 & A_623;
assign w2337 = (~w2336 & w2330) | (~w2336 & w13289) | (w2330 & w13289);
assign w2338 = A_619 & A_620;
assign w2339 = (~w2338 & w2323) | (~w2338 & w13290) | (w2323 & w13290);
assign w2340 = ~w2337 & w2339;
assign w2341 = w2337 & ~w2339;
assign w2342 = ~w2340 & ~w2341;
assign w2343 = ~w2325 & ~w2332;
assign w2344 = ~w2342 & w2343;
assign w2345 = ~w2337 & ~w2339;
assign w2346 = ~w2344 & ~w2345;
assign w2347 = w2343 & w2342;
assign w2348 = ~w2342 & ~w2343;
assign w2349 = ~w2347 & ~w2348;
assign w2350 = ~w2346 & ~w2349;
assign w2351 = ~w2335 & ~w2350;
assign w2352 = ~w2318 & w2351;
assign w2353 = w2318 & ~w2351;
assign w2354 = ~w2352 & ~w2353;
assign w2355 = ~A_613 & A_614;
assign w2356 = A_613 & ~A_614;
assign w2357 = A_615 & ~w2356;
assign w2358 = ~w2355 & w2357;
assign w2359 = ~w2355 & ~w2356;
assign w2360 = ~A_615 & ~w2359;
assign w2361 = ~w2358 & ~w2360;
assign w2362 = ~A_616 & A_617;
assign w2363 = A_616 & ~A_617;
assign w2364 = A_618 & ~w2363;
assign w2365 = ~w2362 & w2364;
assign w2366 = ~w2362 & ~w2363;
assign w2367 = ~A_618 & ~w2366;
assign w2368 = ~w2365 & ~w2367;
assign w2369 = ~w2361 & w2368;
assign w2370 = w2361 & ~w2368;
assign w2371 = ~w2369 & ~w2370;
assign w2372 = A_616 & A_617;
assign w2373 = (~w2372 & w2366) | (~w2372 & w13291) | (w2366 & w13291);
assign w2374 = A_613 & A_614;
assign w2375 = (~w2374 & w2359) | (~w2374 & w13292) | (w2359 & w13292);
assign w2376 = ~w2373 & w2375;
assign w2377 = w2373 & ~w2375;
assign w2378 = ~w2376 & ~w2377;
assign w2379 = ~w2361 & ~w2368;
assign w2380 = ~w2378 & w2379;
assign w2381 = ~w2373 & ~w2375;
assign w2382 = ~w2380 & ~w2381;
assign w2383 = w2379 & w2378;
assign w2384 = ~w2378 & ~w2379;
assign w2385 = ~w2383 & ~w2384;
assign w2386 = ~w2382 & ~w2385;
assign w2387 = ~w2371 & ~w2386;
assign w2388 = ~A_607 & A_608;
assign w2389 = A_607 & ~A_608;
assign w2390 = A_609 & ~w2389;
assign w2391 = ~w2388 & w2390;
assign w2392 = ~w2388 & ~w2389;
assign w2393 = ~A_609 & ~w2392;
assign w2394 = ~w2391 & ~w2393;
assign w2395 = ~A_610 & A_611;
assign w2396 = A_610 & ~A_611;
assign w2397 = A_612 & ~w2396;
assign w2398 = ~w2395 & w2397;
assign w2399 = ~w2395 & ~w2396;
assign w2400 = ~A_612 & ~w2399;
assign w2401 = ~w2398 & ~w2400;
assign w2402 = ~w2394 & w2401;
assign w2403 = w2394 & ~w2401;
assign w2404 = ~w2402 & ~w2403;
assign w2405 = A_610 & A_611;
assign w2406 = (~w2405 & w2399) | (~w2405 & w13293) | (w2399 & w13293);
assign w2407 = A_607 & A_608;
assign w2408 = (~w2407 & w2392) | (~w2407 & w13294) | (w2392 & w13294);
assign w2409 = ~w2406 & w2408;
assign w2410 = w2406 & ~w2408;
assign w2411 = ~w2409 & ~w2410;
assign w2412 = ~w2394 & ~w2401;
assign w2413 = ~w2411 & w2412;
assign w2414 = ~w2406 & ~w2408;
assign w2415 = ~w2413 & ~w2414;
assign w2416 = w2412 & w2411;
assign w2417 = ~w2411 & ~w2412;
assign w2418 = ~w2416 & ~w2417;
assign w2419 = ~w2415 & ~w2418;
assign w2420 = ~w2404 & ~w2419;
assign w2421 = ~w2387 & w2420;
assign w2422 = w2387 & ~w2420;
assign w2423 = ~w2421 & ~w2422;
assign w2424 = ~w2354 & w2423;
assign w2425 = w2354 & ~w2423;
assign w2426 = ~w2424 & ~w2425;
assign w2427 = ~w2285 & w2426;
assign w2428 = w2285 & ~w2426;
assign w2429 = ~w2427 & ~w2428;
assign w2430 = ~A_601 & A_602;
assign w2431 = A_601 & ~A_602;
assign w2432 = A_603 & ~w2431;
assign w2433 = ~w2430 & w2432;
assign w2434 = ~w2430 & ~w2431;
assign w2435 = ~A_603 & ~w2434;
assign w2436 = ~w2433 & ~w2435;
assign w2437 = ~A_604 & A_605;
assign w2438 = A_604 & ~A_605;
assign w2439 = A_606 & ~w2438;
assign w2440 = ~w2437 & w2439;
assign w2441 = ~w2437 & ~w2438;
assign w2442 = ~A_606 & ~w2441;
assign w2443 = ~w2440 & ~w2442;
assign w2444 = ~w2436 & w2443;
assign w2445 = w2436 & ~w2443;
assign w2446 = ~w2444 & ~w2445;
assign w2447 = A_604 & A_605;
assign w2448 = (~w2447 & w2441) | (~w2447 & w13295) | (w2441 & w13295);
assign w2449 = A_601 & A_602;
assign w2450 = (~w2449 & w2434) | (~w2449 & w13296) | (w2434 & w13296);
assign w2451 = ~w2448 & w2450;
assign w2452 = w2448 & ~w2450;
assign w2453 = ~w2451 & ~w2452;
assign w2454 = ~w2436 & ~w2443;
assign w2455 = ~w2453 & w2454;
assign w2456 = ~w2448 & ~w2450;
assign w2457 = ~w2455 & ~w2456;
assign w2458 = w2454 & w2453;
assign w2459 = ~w2453 & ~w2454;
assign w2460 = ~w2458 & ~w2459;
assign w2461 = ~w2457 & ~w2460;
assign w2462 = ~w2446 & ~w2461;
assign w2463 = ~A_595 & A_596;
assign w2464 = A_595 & ~A_596;
assign w2465 = A_597 & ~w2464;
assign w2466 = ~w2463 & w2465;
assign w2467 = ~w2463 & ~w2464;
assign w2468 = ~A_597 & ~w2467;
assign w2469 = ~w2466 & ~w2468;
assign w2470 = ~A_598 & A_599;
assign w2471 = A_598 & ~A_599;
assign w2472 = A_600 & ~w2471;
assign w2473 = ~w2470 & w2472;
assign w2474 = ~w2470 & ~w2471;
assign w2475 = ~A_600 & ~w2474;
assign w2476 = ~w2473 & ~w2475;
assign w2477 = ~w2469 & w2476;
assign w2478 = w2469 & ~w2476;
assign w2479 = ~w2477 & ~w2478;
assign w2480 = A_598 & A_599;
assign w2481 = (~w2480 & w2474) | (~w2480 & w13297) | (w2474 & w13297);
assign w2482 = A_595 & A_596;
assign w2483 = (~w2482 & w2467) | (~w2482 & w13298) | (w2467 & w13298);
assign w2484 = ~w2481 & w2483;
assign w2485 = w2481 & ~w2483;
assign w2486 = ~w2484 & ~w2485;
assign w2487 = ~w2469 & ~w2476;
assign w2488 = ~w2486 & w2487;
assign w2489 = ~w2481 & ~w2483;
assign w2490 = ~w2488 & ~w2489;
assign w2491 = w2487 & w2486;
assign w2492 = ~w2486 & ~w2487;
assign w2493 = ~w2491 & ~w2492;
assign w2494 = ~w2490 & ~w2493;
assign w2495 = ~w2479 & ~w2494;
assign w2496 = ~w2462 & w2495;
assign w2497 = w2462 & ~w2495;
assign w2498 = ~w2496 & ~w2497;
assign w2499 = ~A_589 & A_590;
assign w2500 = A_589 & ~A_590;
assign w2501 = A_591 & ~w2500;
assign w2502 = ~w2499 & w2501;
assign w2503 = ~w2499 & ~w2500;
assign w2504 = ~A_591 & ~w2503;
assign w2505 = ~w2502 & ~w2504;
assign w2506 = ~A_592 & A_593;
assign w2507 = A_592 & ~A_593;
assign w2508 = A_594 & ~w2507;
assign w2509 = ~w2506 & w2508;
assign w2510 = ~w2506 & ~w2507;
assign w2511 = ~A_594 & ~w2510;
assign w2512 = ~w2509 & ~w2511;
assign w2513 = ~w2505 & w2512;
assign w2514 = w2505 & ~w2512;
assign w2515 = ~w2513 & ~w2514;
assign w2516 = A_592 & A_593;
assign w2517 = (~w2516 & w2510) | (~w2516 & w13299) | (w2510 & w13299);
assign w2518 = A_589 & A_590;
assign w2519 = (~w2518 & w2503) | (~w2518 & w13300) | (w2503 & w13300);
assign w2520 = ~w2517 & w2519;
assign w2521 = w2517 & ~w2519;
assign w2522 = ~w2520 & ~w2521;
assign w2523 = ~w2505 & ~w2512;
assign w2524 = ~w2522 & w2523;
assign w2525 = ~w2517 & ~w2519;
assign w2526 = ~w2524 & ~w2525;
assign w2527 = w2523 & w2522;
assign w2528 = ~w2522 & ~w2523;
assign w2529 = ~w2527 & ~w2528;
assign w2530 = ~w2526 & ~w2529;
assign w2531 = ~w2515 & ~w2530;
assign w2532 = ~A_583 & A_584;
assign w2533 = A_583 & ~A_584;
assign w2534 = A_585 & ~w2533;
assign w2535 = ~w2532 & w2534;
assign w2536 = ~w2532 & ~w2533;
assign w2537 = ~A_585 & ~w2536;
assign w2538 = ~w2535 & ~w2537;
assign w2539 = ~A_586 & A_587;
assign w2540 = A_586 & ~A_587;
assign w2541 = A_588 & ~w2540;
assign w2542 = ~w2539 & w2541;
assign w2543 = ~w2539 & ~w2540;
assign w2544 = ~A_588 & ~w2543;
assign w2545 = ~w2542 & ~w2544;
assign w2546 = ~w2538 & w2545;
assign w2547 = w2538 & ~w2545;
assign w2548 = ~w2546 & ~w2547;
assign w2549 = A_586 & A_587;
assign w2550 = (~w2549 & w2543) | (~w2549 & w13301) | (w2543 & w13301);
assign w2551 = A_583 & A_584;
assign w2552 = (~w2551 & w2536) | (~w2551 & w13302) | (w2536 & w13302);
assign w2553 = ~w2550 & w2552;
assign w2554 = w2550 & ~w2552;
assign w2555 = ~w2553 & ~w2554;
assign w2556 = ~w2538 & ~w2545;
assign w2557 = ~w2555 & w2556;
assign w2558 = ~w2550 & ~w2552;
assign w2559 = ~w2557 & ~w2558;
assign w2560 = w2556 & w2555;
assign w2561 = ~w2555 & ~w2556;
assign w2562 = ~w2560 & ~w2561;
assign w2563 = ~w2559 & ~w2562;
assign w2564 = ~w2548 & ~w2563;
assign w2565 = ~w2531 & w2564;
assign w2566 = w2531 & ~w2564;
assign w2567 = ~w2565 & ~w2566;
assign w2568 = ~w2498 & w2567;
assign w2569 = w2498 & ~w2567;
assign w2570 = ~w2568 & ~w2569;
assign w2571 = ~A_577 & A_578;
assign w2572 = A_577 & ~A_578;
assign w2573 = A_579 & ~w2572;
assign w2574 = ~w2571 & w2573;
assign w2575 = ~w2571 & ~w2572;
assign w2576 = ~A_579 & ~w2575;
assign w2577 = ~w2574 & ~w2576;
assign w2578 = ~A_580 & A_581;
assign w2579 = A_580 & ~A_581;
assign w2580 = A_582 & ~w2579;
assign w2581 = ~w2578 & w2580;
assign w2582 = ~w2578 & ~w2579;
assign w2583 = ~A_582 & ~w2582;
assign w2584 = ~w2581 & ~w2583;
assign w2585 = ~w2577 & w2584;
assign w2586 = w2577 & ~w2584;
assign w2587 = ~w2585 & ~w2586;
assign w2588 = A_580 & A_581;
assign w2589 = (~w2588 & w2582) | (~w2588 & w13303) | (w2582 & w13303);
assign w2590 = A_577 & A_578;
assign w2591 = (~w2590 & w2575) | (~w2590 & w13304) | (w2575 & w13304);
assign w2592 = ~w2589 & w2591;
assign w2593 = w2589 & ~w2591;
assign w2594 = ~w2592 & ~w2593;
assign w2595 = ~w2577 & ~w2584;
assign w2596 = ~w2594 & w2595;
assign w2597 = ~w2589 & ~w2591;
assign w2598 = ~w2596 & ~w2597;
assign w2599 = w2595 & w2594;
assign w2600 = ~w2594 & ~w2595;
assign w2601 = ~w2599 & ~w2600;
assign w2602 = ~w2598 & ~w2601;
assign w2603 = ~w2587 & ~w2602;
assign w2604 = ~A_571 & A_572;
assign w2605 = A_571 & ~A_572;
assign w2606 = A_573 & ~w2605;
assign w2607 = ~w2604 & w2606;
assign w2608 = ~w2604 & ~w2605;
assign w2609 = ~A_573 & ~w2608;
assign w2610 = ~w2607 & ~w2609;
assign w2611 = ~A_574 & A_575;
assign w2612 = A_574 & ~A_575;
assign w2613 = A_576 & ~w2612;
assign w2614 = ~w2611 & w2613;
assign w2615 = ~w2611 & ~w2612;
assign w2616 = ~A_576 & ~w2615;
assign w2617 = ~w2614 & ~w2616;
assign w2618 = ~w2610 & w2617;
assign w2619 = w2610 & ~w2617;
assign w2620 = ~w2618 & ~w2619;
assign w2621 = A_574 & A_575;
assign w2622 = (~w2621 & w2615) | (~w2621 & w13305) | (w2615 & w13305);
assign w2623 = A_571 & A_572;
assign w2624 = (~w2623 & w2608) | (~w2623 & w13306) | (w2608 & w13306);
assign w2625 = ~w2622 & w2624;
assign w2626 = w2622 & ~w2624;
assign w2627 = ~w2625 & ~w2626;
assign w2628 = ~w2610 & ~w2617;
assign w2629 = ~w2627 & w2628;
assign w2630 = ~w2622 & ~w2624;
assign w2631 = ~w2629 & ~w2630;
assign w2632 = w2628 & w2627;
assign w2633 = ~w2627 & ~w2628;
assign w2634 = ~w2632 & ~w2633;
assign w2635 = ~w2631 & ~w2634;
assign w2636 = ~w2620 & ~w2635;
assign w2637 = ~w2603 & w2636;
assign w2638 = w2603 & ~w2636;
assign w2639 = ~w2637 & ~w2638;
assign w2640 = ~A_565 & A_566;
assign w2641 = A_565 & ~A_566;
assign w2642 = A_567 & ~w2641;
assign w2643 = ~w2640 & w2642;
assign w2644 = ~w2640 & ~w2641;
assign w2645 = ~A_567 & ~w2644;
assign w2646 = ~w2643 & ~w2645;
assign w2647 = ~A_568 & A_569;
assign w2648 = A_568 & ~A_569;
assign w2649 = A_570 & ~w2648;
assign w2650 = ~w2647 & w2649;
assign w2651 = ~w2647 & ~w2648;
assign w2652 = ~A_570 & ~w2651;
assign w2653 = ~w2650 & ~w2652;
assign w2654 = ~w2646 & w2653;
assign w2655 = w2646 & ~w2653;
assign w2656 = ~w2654 & ~w2655;
assign w2657 = A_568 & A_569;
assign w2658 = (~w2657 & w2651) | (~w2657 & w13307) | (w2651 & w13307);
assign w2659 = A_565 & A_566;
assign w2660 = (~w2659 & w2644) | (~w2659 & w13308) | (w2644 & w13308);
assign w2661 = ~w2658 & w2660;
assign w2662 = w2658 & ~w2660;
assign w2663 = ~w2661 & ~w2662;
assign w2664 = ~w2646 & ~w2653;
assign w2665 = ~w2663 & w2664;
assign w2666 = ~w2658 & ~w2660;
assign w2667 = ~w2665 & ~w2666;
assign w2668 = w2664 & w2663;
assign w2669 = ~w2663 & ~w2664;
assign w2670 = ~w2668 & ~w2669;
assign w2671 = ~w2667 & ~w2670;
assign w2672 = ~w2656 & ~w2671;
assign w2673 = ~A_559 & A_560;
assign w2674 = A_559 & ~A_560;
assign w2675 = A_561 & ~w2674;
assign w2676 = ~w2673 & w2675;
assign w2677 = ~w2673 & ~w2674;
assign w2678 = ~A_561 & ~w2677;
assign w2679 = ~w2676 & ~w2678;
assign w2680 = ~A_562 & A_563;
assign w2681 = A_562 & ~A_563;
assign w2682 = A_564 & ~w2681;
assign w2683 = ~w2680 & w2682;
assign w2684 = ~w2680 & ~w2681;
assign w2685 = ~A_564 & ~w2684;
assign w2686 = ~w2683 & ~w2685;
assign w2687 = ~w2679 & w2686;
assign w2688 = w2679 & ~w2686;
assign w2689 = ~w2687 & ~w2688;
assign w2690 = A_562 & A_563;
assign w2691 = (~w2690 & w2684) | (~w2690 & w13309) | (w2684 & w13309);
assign w2692 = A_559 & A_560;
assign w2693 = (~w2692 & w2677) | (~w2692 & w13310) | (w2677 & w13310);
assign w2694 = ~w2691 & w2693;
assign w2695 = w2691 & ~w2693;
assign w2696 = ~w2694 & ~w2695;
assign w2697 = ~w2679 & ~w2686;
assign w2698 = ~w2696 & w2697;
assign w2699 = ~w2691 & ~w2693;
assign w2700 = ~w2698 & ~w2699;
assign w2701 = w2697 & w2696;
assign w2702 = ~w2696 & ~w2697;
assign w2703 = ~w2701 & ~w2702;
assign w2704 = ~w2700 & ~w2703;
assign w2705 = ~w2689 & ~w2704;
assign w2706 = ~w2672 & w2705;
assign w2707 = w2672 & ~w2705;
assign w2708 = ~w2706 & ~w2707;
assign w2709 = ~w2639 & w2708;
assign w2710 = w2639 & ~w2708;
assign w2711 = ~w2709 & ~w2710;
assign w2712 = ~w2570 & w2711;
assign w2713 = w2570 & ~w2711;
assign w2714 = ~w2712 & ~w2713;
assign w2715 = ~w2429 & w2714;
assign w2716 = w2429 & ~w2714;
assign w2717 = ~w2715 & ~w2716;
assign w2718 = ~w2144 & w2717;
assign w2719 = w2144 & ~w2717;
assign w2720 = ~w2718 & ~w2719;
assign w2721 = ~w1557 & w1560;
assign w2722 = w1557 & ~w1560;
assign w2723 = ~w2721 & ~w2722;
assign w2724 = ~w2720 & ~w2723;
assign w2725 = (w2724 & w1570) | (w2724 & w13813) | (w1570 & w13813);
assign w2726 = ~w1566 & w2725;
assign w2727 = (~w2724 & w1571) | (~w2724 & w13814) | (w1571 & w13814);
assign w2728 = ~w2726 & ~w2727;
assign w2729 = ~w2548 & ~w2559;
assign w2730 = ~w2562 & ~w2729;
assign w2731 = ~w2515 & ~w2548;
assign w2732 = ~w2530 & w2731;
assign w2733 = ~w2563 & w2732;
assign w2734 = ~w2515 & ~w2526;
assign w2735 = ~w2529 & ~w2734;
assign w2736 = ~w2733 & w2735;
assign w2737 = w2733 & ~w2735;
assign w2738 = ~w2736 & ~w2737;
assign w2739 = ~w2730 & ~w2738;
assign w2740 = ~w2733 & ~w2735;
assign w2741 = ~w2529 & w2731;
assign w2742 = ~w2530 & w2741;
assign w2743 = ~w2563 & ~w2734;
assign w2744 = w2742 & w2743;
assign w2745 = (w2730 & w2740) | (w2730 & w13689) | (w2740 & w13689);
assign w2746 = ~w2739 & ~w2745;
assign w2747 = ~w2479 & ~w2490;
assign w2748 = ~w2493 & ~w2747;
assign w2749 = ~w2446 & ~w2479;
assign w2750 = ~w2461 & w2749;
assign w2751 = ~w2494 & w2750;
assign w2752 = ~w2446 & ~w2457;
assign w2753 = ~w2460 & ~w2752;
assign w2754 = ~w2751 & ~w2753;
assign w2755 = ~w2460 & w2749;
assign w2756 = ~w2461 & w2755;
assign w2757 = ~w2494 & ~w2752;
assign w2758 = w2756 & w2757;
assign w2759 = (w2748 & w2754) | (w2748 & w13496) | (w2754 & w13496);
assign w2760 = ~w2751 & w2753;
assign w2761 = w2751 & ~w2753;
assign w2762 = ~w2760 & ~w2761;
assign w2763 = ~w2748 & ~w2762;
assign w2764 = ~w2498 & ~w2567;
assign w2765 = ~w2763 & w13497;
assign w2766 = (w2764 & w2763) | (w2764 & w13690) | (w2763 & w13690);
assign w2767 = ~w2765 & ~w2766;
assign w2768 = ~w2746 & ~w2767;
assign w2769 = ~w2763 & w13498;
assign w2770 = (~w2764 & w2763) | (~w2764 & w13691) | (w2763 & w13691);
assign w2771 = (w2746 & w2770) | (w2746 & w13499) | (w2770 & w13499);
assign w2772 = ~w2570 & ~w2711;
assign w2773 = w2772 & ~w2771;
assign w2774 = ~w2768 & w2773;
assign w2775 = ~w2768 & ~w2771;
assign w2776 = ~w2772 & ~w2775;
assign w2777 = ~w2620 & ~w2631;
assign w2778 = ~w2634 & ~w2777;
assign w2779 = ~w2587 & ~w2620;
assign w2780 = ~w2602 & w2779;
assign w2781 = ~w2635 & w2780;
assign w2782 = ~w2587 & ~w2598;
assign w2783 = ~w2601 & ~w2782;
assign w2784 = ~w2781 & ~w2783;
assign w2785 = ~w2601 & w2779;
assign w2786 = ~w2602 & w2785;
assign w2787 = ~w2635 & ~w2782;
assign w2788 = w2786 & w2787;
assign w2789 = (w2778 & w2784) | (w2778 & w13692) | (w2784 & w13692);
assign w2790 = ~w2781 & w2783;
assign w2791 = w2781 & ~w2783;
assign w2792 = ~w2790 & ~w2791;
assign w2793 = ~w2778 & ~w2792;
assign w2794 = ~w2639 & ~w2708;
assign w2795 = ~w2793 & w13693;
assign w2796 = (~w2794 & w2793) | (~w2794 & w13694) | (w2793 & w13694);
assign w2797 = ~w2795 & ~w2796;
assign w2798 = ~w2689 & ~w2700;
assign w2799 = ~w2703 & ~w2798;
assign w2800 = ~w2656 & ~w2689;
assign w2801 = ~w2671 & w2800;
assign w2802 = ~w2704 & w2801;
assign w2803 = ~w2656 & ~w2667;
assign w2804 = ~w2670 & ~w2803;
assign w2805 = ~w2802 & w2804;
assign w2806 = w2802 & ~w2804;
assign w2807 = ~w2805 & ~w2806;
assign w2808 = ~w2799 & ~w2807;
assign w2809 = ~w2802 & ~w2804;
assign w2810 = ~w2670 & w2800;
assign w2811 = ~w2671 & w2810;
assign w2812 = ~w2704 & ~w2803;
assign w2813 = w2811 & w2812;
assign w2814 = (w2799 & w2809) | (w2799 & w13815) | (w2809 & w13815);
assign w2815 = ~w2808 & ~w2814;
assign w2816 = ~w2797 & w2815;
assign w2817 = ~w2793 & w13695;
assign w2818 = (w2794 & w2793) | (w2794 & w13816) | (w2793 & w13816);
assign w2819 = (~w2815 & w2818) | (~w2815 & w13696) | (w2818 & w13696);
assign w2820 = ~w2816 & ~w2819;
assign w2821 = (w2820 & w2776) | (w2820 & w13817) | (w2776 & w13817);
assign w2822 = ~w2772 & ~w2771;
assign w2823 = ~w2768 & w2822;
assign w2824 = w2772 & ~w2775;
assign w2825 = (~w2820 & w2824) | (~w2820 & w13818) | (w2824 & w13818);
assign w2826 = ~w2821 & ~w2825;
assign w2827 = ~w2335 & ~w2346;
assign w2828 = ~w2349 & ~w2827;
assign w2829 = ~w2302 & ~w2335;
assign w2830 = ~w2317 & w2829;
assign w2831 = ~w2350 & w2830;
assign w2832 = ~w2302 & ~w2313;
assign w2833 = ~w2316 & ~w2832;
assign w2834 = ~w2831 & ~w2833;
assign w2835 = ~w2316 & w2829;
assign w2836 = ~w2317 & w2835;
assign w2837 = ~w2350 & ~w2832;
assign w2838 = w2836 & w2837;
assign w2839 = (w2828 & w2834) | (w2828 & w13697) | (w2834 & w13697);
assign w2840 = ~w2831 & w2833;
assign w2841 = w2831 & ~w2833;
assign w2842 = ~w2840 & ~w2841;
assign w2843 = ~w2828 & ~w2842;
assign w2844 = ~w2354 & ~w2423;
assign w2845 = ~w2843 & w13698;
assign w2846 = (~w2844 & w2843) | (~w2844 & w13699) | (w2843 & w13699);
assign w2847 = ~w2845 & ~w2846;
assign w2848 = ~w2404 & ~w2415;
assign w2849 = ~w2418 & ~w2848;
assign w2850 = ~w2371 & ~w2404;
assign w2851 = ~w2386 & w2850;
assign w2852 = ~w2419 & w2851;
assign w2853 = ~w2371 & ~w2382;
assign w2854 = ~w2385 & ~w2853;
assign w2855 = ~w2852 & w2854;
assign w2856 = w2852 & ~w2854;
assign w2857 = ~w2855 & ~w2856;
assign w2858 = ~w2849 & ~w2857;
assign w2859 = ~w2852 & ~w2854;
assign w2860 = ~w2385 & w2850;
assign w2861 = ~w2386 & w2860;
assign w2862 = ~w2419 & ~w2853;
assign w2863 = w2861 & w2862;
assign w2864 = (w2849 & w2859) | (w2849 & w13819) | (w2859 & w13819);
assign w2865 = ~w2858 & ~w2864;
assign w2866 = ~w2847 & w2865;
assign w2867 = ~w2843 & w13700;
assign w2868 = (w2844 & w2843) | (w2844 & w13820) | (w2843 & w13820);
assign w2869 = (~w2865 & w2868) | (~w2865 & w13701) | (w2868 & w13701);
assign w2870 = ~w2866 & ~w2869;
assign w2871 = ~w2263 & ~w2274;
assign w2872 = ~w2277 & ~w2871;
assign w2873 = ~w2230 & ~w2263;
assign w2874 = ~w2245 & w2873;
assign w2875 = ~w2278 & w2874;
assign w2876 = ~w2230 & ~w2241;
assign w2877 = ~w2244 & ~w2876;
assign w2878 = ~w2875 & w2877;
assign w2879 = w2875 & ~w2877;
assign w2880 = ~w2878 & ~w2879;
assign w2881 = ~w2872 & ~w2880;
assign w2882 = ~w2875 & ~w2877;
assign w2883 = ~w2244 & w2873;
assign w2884 = ~w2245 & w2883;
assign w2885 = ~w2278 & ~w2876;
assign w2886 = w2884 & w2885;
assign w2887 = (w2872 & w2882) | (w2872 & w13702) | (w2882 & w13702);
assign w2888 = ~w2881 & ~w2887;
assign w2889 = ~w2194 & ~w2205;
assign w2890 = ~w2208 & ~w2889;
assign w2891 = ~w2161 & ~w2194;
assign w2892 = ~w2176 & w2891;
assign w2893 = ~w2209 & w2892;
assign w2894 = ~w2161 & ~w2172;
assign w2895 = ~w2175 & ~w2894;
assign w2896 = ~w2893 & ~w2895;
assign w2897 = ~w2175 & w2891;
assign w2898 = ~w2176 & w2897;
assign w2899 = ~w2209 & ~w2894;
assign w2900 = w2898 & w2899;
assign w2901 = (w2890 & w2896) | (w2890 & w13500) | (w2896 & w13500);
assign w2902 = ~w2893 & w2895;
assign w2903 = w2893 & ~w2895;
assign w2904 = ~w2902 & ~w2903;
assign w2905 = ~w2890 & ~w2904;
assign w2906 = ~w2213 & ~w2282;
assign w2907 = ~w2905 & w13501;
assign w2908 = (w2906 & w2905) | (w2906 & w13502) | (w2905 & w13502);
assign w2909 = ~w2907 & ~w2908;
assign w2910 = ~w2888 & ~w2909;
assign w2911 = ~w2905 & w13503;
assign w2912 = (~w2906 & w2905) | (~w2906 & w13703) | (w2905 & w13703);
assign w2913 = (w2888 & w2912) | (w2888 & w13504) | (w2912 & w13504);
assign w2914 = ~w2285 & ~w2426;
assign w2915 = ~w2914 & ~w2913;
assign w2916 = ~w2910 & w2915;
assign w2917 = ~w2910 & ~w2913;
assign w2918 = w2914 & ~w2917;
assign w2919 = (~w2870 & w2918) | (~w2870 & w13704) | (w2918 & w13704);
assign w2920 = w2914 & ~w2913;
assign w2921 = ~w2910 & w2920;
assign w2922 = ~w2914 & ~w2917;
assign w2923 = ~w2921 & ~w2922;
assign w2924 = (w2870 & w2922) | (w2870 & w13821) | (w2922 & w13821);
assign w2925 = ~w2429 & ~w2714;
assign w2926 = (~w2925 & w2923) | (~w2925 & w13705) | (w2923 & w13705);
assign w2927 = ~w2919 & w2926;
assign w2928 = ~w2919 & ~w2924;
assign w2929 = w2925 & ~w2928;
assign w2930 = ~w2927 & ~w2929;
assign w2931 = ~w2826 & ~w2930;
assign w2932 = (w2925 & w2923) | (w2925 & w13706) | (w2923 & w13706);
assign w2933 = ~w2919 & w2932;
assign w2934 = (~w2925 & w2924) | (~w2925 & w13707) | (w2924 & w13707);
assign w2935 = ~w2933 & ~w2934;
assign w2936 = w2826 & ~w2935;
assign w2937 = ~w2144 & ~w2717;
assign w2938 = (w2937 & w2935) | (w2937 & w13822) | (w2935 & w13822);
assign w2939 = ~w2931 & w2938;
assign w2940 = ~w2931 & ~w2936;
assign w2941 = ~w2937 & ~w2940;
assign w2942 = ~w2047 & ~w2058;
assign w2943 = ~w2061 & ~w2942;
assign w2944 = ~w2014 & ~w2047;
assign w2945 = ~w2029 & w2944;
assign w2946 = ~w2062 & w2945;
assign w2947 = ~w2014 & ~w2025;
assign w2948 = ~w2028 & ~w2947;
assign w2949 = ~w2946 & ~w2948;
assign w2950 = ~w2028 & w2944;
assign w2951 = ~w2029 & w2950;
assign w2952 = ~w2062 & ~w2947;
assign w2953 = w2951 & w2952;
assign w2954 = (w2943 & w2949) | (w2943 & w13708) | (w2949 & w13708);
assign w2955 = ~w2946 & w2948;
assign w2956 = w2946 & ~w2948;
assign w2957 = ~w2955 & ~w2956;
assign w2958 = ~w2943 & ~w2957;
assign w2959 = ~w2066 & ~w2135;
assign w2960 = ~w2958 & w13709;
assign w2961 = (~w2959 & w2958) | (~w2959 & w13710) | (w2958 & w13710);
assign w2962 = ~w2960 & ~w2961;
assign w2963 = ~w2116 & ~w2127;
assign w2964 = ~w2130 & ~w2963;
assign w2965 = ~w2083 & ~w2116;
assign w2966 = ~w2098 & w2965;
assign w2967 = ~w2131 & w2966;
assign w2968 = ~w2083 & ~w2094;
assign w2969 = ~w2097 & ~w2968;
assign w2970 = ~w2967 & w2969;
assign w2971 = w2967 & ~w2969;
assign w2972 = ~w2970 & ~w2971;
assign w2973 = ~w2964 & ~w2972;
assign w2974 = ~w2967 & ~w2969;
assign w2975 = ~w2097 & w2965;
assign w2976 = ~w2098 & w2975;
assign w2977 = ~w2131 & ~w2968;
assign w2978 = w2976 & w2977;
assign w2979 = (w2964 & w2974) | (w2964 & w13823) | (w2974 & w13823);
assign w2980 = ~w2973 & ~w2979;
assign w2981 = ~w2962 & w2980;
assign w2982 = ~w2958 & w13711;
assign w2983 = (w2959 & w2958) | (w2959 & w13824) | (w2958 & w13824);
assign w2984 = (~w2980 & w2983) | (~w2980 & w13712) | (w2983 & w13712);
assign w2985 = ~w2981 & ~w2984;
assign w2986 = ~w1975 & ~w1986;
assign w2987 = ~w1989 & ~w2986;
assign w2988 = ~w1942 & ~w1975;
assign w2989 = ~w1957 & w2988;
assign w2990 = ~w1990 & w2989;
assign w2991 = ~w1942 & ~w1953;
assign w2992 = ~w1956 & ~w2991;
assign w2993 = ~w2990 & w2992;
assign w2994 = w2990 & ~w2992;
assign w2995 = ~w2993 & ~w2994;
assign w2996 = ~w2987 & ~w2995;
assign w2997 = ~w2990 & ~w2992;
assign w2998 = ~w1956 & w2988;
assign w2999 = ~w1957 & w2998;
assign w3000 = ~w1990 & ~w2991;
assign w3001 = w2999 & w3000;
assign w3002 = (w2987 & w2997) | (w2987 & w13713) | (w2997 & w13713);
assign w3003 = ~w2996 & ~w3002;
assign w3004 = ~w1906 & ~w1917;
assign w3005 = ~w1920 & ~w3004;
assign w3006 = ~w1873 & ~w1906;
assign w3007 = ~w1888 & w3006;
assign w3008 = ~w1921 & w3007;
assign w3009 = ~w1873 & ~w1884;
assign w3010 = ~w1887 & ~w3009;
assign w3011 = ~w3008 & ~w3010;
assign w3012 = ~w1887 & w3006;
assign w3013 = ~w1888 & w3012;
assign w3014 = ~w1921 & ~w3009;
assign w3015 = w3013 & w3014;
assign w3016 = (w3005 & w3011) | (w3005 & w13505) | (w3011 & w13505);
assign w3017 = ~w3008 & w3010;
assign w3018 = w3008 & ~w3010;
assign w3019 = ~w3017 & ~w3018;
assign w3020 = ~w3005 & ~w3019;
assign w3021 = ~w1925 & ~w1994;
assign w3022 = ~w3020 & w13506;
assign w3023 = (w3021 & w3020) | (w3021 & w13507) | (w3020 & w13507);
assign w3024 = ~w3022 & ~w3023;
assign w3025 = ~w3003 & ~w3024;
assign w3026 = ~w3020 & w13508;
assign w3027 = (~w3021 & w3020) | (~w3021 & w13714) | (w3020 & w13714);
assign w3028 = (w3003 & w3027) | (w3003 & w13509) | (w3027 & w13509);
assign w3029 = ~w1997 & ~w2138;
assign w3030 = ~w3029 & ~w3028;
assign w3031 = ~w3025 & w3030;
assign w3032 = ~w3025 & ~w3028;
assign w3033 = w3029 & ~w3032;
assign w3034 = (~w2985 & w3033) | (~w2985 & w13825) | (w3033 & w13825);
assign w3035 = w3029 & ~w3028;
assign w3036 = ~w3025 & w3035;
assign w3037 = ~w3029 & ~w3032;
assign w3038 = (w2985 & w3037) | (w2985 & w13715) | (w3037 & w13715);
assign w3039 = ~w1856 & ~w2141;
assign w3040 = ~w3038 & w3039;
assign w3041 = ~w3034 & w3040;
assign w3042 = ~w3034 & ~w3038;
assign w3043 = ~w3039 & ~w3042;
assign w3044 = ~w3041 & ~w3043;
assign w3045 = ~w1831 & ~w1842;
assign w3046 = ~w1845 & ~w3045;
assign w3047 = ~w1798 & ~w1831;
assign w3048 = ~w1813 & w3047;
assign w3049 = ~w1846 & w3048;
assign w3050 = ~w1798 & ~w1809;
assign w3051 = ~w1812 & ~w3050;
assign w3052 = ~w3049 & w3051;
assign w3053 = w3049 & ~w3051;
assign w3054 = ~w3052 & ~w3053;
assign w3055 = ~w3046 & ~w3054;
assign w3056 = ~w3049 & ~w3051;
assign w3057 = ~w1812 & w3047;
assign w3058 = ~w1813 & w3057;
assign w3059 = ~w1846 & ~w3050;
assign w3060 = w3058 & w3059;
assign w3061 = (w3046 & w3056) | (w3046 & w13716) | (w3056 & w13716);
assign w3062 = ~w3055 & ~w3061;
assign w3063 = ~w1762 & ~w1773;
assign w3064 = ~w1776 & ~w3063;
assign w3065 = ~w1729 & ~w1762;
assign w3066 = ~w1744 & w3065;
assign w3067 = ~w1777 & w3066;
assign w3068 = ~w1729 & ~w1740;
assign w3069 = ~w1743 & ~w3068;
assign w3070 = ~w3067 & ~w3069;
assign w3071 = ~w1743 & w3065;
assign w3072 = ~w1744 & w3071;
assign w3073 = ~w1777 & ~w3068;
assign w3074 = w3072 & w3073;
assign w3075 = (w3064 & w3070) | (w3064 & w13510) | (w3070 & w13510);
assign w3076 = ~w3067 & w3069;
assign w3077 = w3067 & ~w3069;
assign w3078 = ~w3076 & ~w3077;
assign w3079 = ~w3064 & ~w3078;
assign w3080 = ~w1781 & ~w1850;
assign w3081 = ~w3079 & w13511;
assign w3082 = (w3080 & w3079) | (w3080 & w13717) | (w3079 & w13717);
assign w3083 = ~w3081 & ~w3082;
assign w3084 = ~w3062 & ~w3083;
assign w3085 = ~w3079 & w13512;
assign w3086 = (~w3080 & w3079) | (~w3080 & w13718) | (w3079 & w13718);
assign w3087 = (w3062 & w3086) | (w3062 & w13513) | (w3086 & w13513);
assign w3088 = ~w1712 & ~w1853;
assign w3089 = w3088 & ~w3087;
assign w3090 = ~w3084 & w3089;
assign w3091 = ~w3084 & ~w3087;
assign w3092 = ~w3088 & ~w3091;
assign w3093 = ~w1690 & ~w1701;
assign w3094 = ~w1704 & ~w3093;
assign w3095 = ~w1657 & ~w1690;
assign w3096 = ~w1672 & w3095;
assign w3097 = ~w1705 & w3096;
assign w3098 = ~w1657 & ~w1668;
assign w3099 = ~w1671 & ~w3098;
assign w3100 = ~w3097 & ~w3099;
assign w3101 = ~w1671 & w3095;
assign w3102 = ~w1672 & w3101;
assign w3103 = ~w1705 & ~w3098;
assign w3104 = w3102 & w3103;
assign w3105 = (w3094 & w3100) | (w3094 & w13719) | (w3100 & w13719);
assign w3106 = ~w3097 & w3099;
assign w3107 = w3097 & ~w3099;
assign w3108 = ~w3106 & ~w3107;
assign w3109 = ~w3094 & ~w3108;
assign w3110 = ~w1640 & ~w1709;
assign w3111 = ~w3109 & w13720;
assign w3112 = (~w3110 & w3109) | (~w3110 & w13721) | (w3109 & w13721);
assign w3113 = ~w3111 & ~w3112;
assign w3114 = ~w1621 & ~w1635;
assign w3115 = ~w1632 & ~w3114;
assign w3116 = ~w1588 & ~w1621;
assign w3117 = ~w1603 & w3116;
assign w3118 = ~w1636 & w3117;
assign w3119 = ~w1588 & ~w1599;
assign w3120 = ~w1602 & ~w3119;
assign w3121 = ~w3118 & w3120;
assign w3122 = w3118 & ~w3120;
assign w3123 = ~w3121 & ~w3122;
assign w3124 = ~w3115 & ~w3123;
assign w3125 = ~w3118 & ~w3120;
assign w3126 = ~w1602 & w3116;
assign w3127 = ~w1603 & w3126;
assign w3128 = ~w1636 & ~w3119;
assign w3129 = w3127 & w3128;
assign w3130 = (w3115 & w3125) | (w3115 & w13826) | (w3125 & w13826);
assign w3131 = ~w3124 & ~w3130;
assign w3132 = ~w3113 & w3131;
assign w3133 = ~w3109 & w13722;
assign w3134 = (w3110 & w3109) | (w3110 & w13827) | (w3109 & w13827);
assign w3135 = (~w3131 & w3134) | (~w3131 & w13723) | (w3134 & w13723);
assign w3136 = ~w3132 & ~w3135;
assign w3137 = (w3136 & w3092) | (w3136 & w13828) | (w3092 & w13828);
assign w3138 = ~w3088 & ~w3087;
assign w3139 = ~w3084 & w3138;
assign w3140 = w3088 & ~w3091;
assign w3141 = (~w3136 & w3140) | (~w3136 & w13829) | (w3140 & w13829);
assign w3142 = ~w3137 & ~w3141;
assign w3143 = ~w3044 & w3142;
assign w3144 = ~w3038 & ~w3039;
assign w3145 = ~w3034 & w3144;
assign w3146 = w3039 & ~w3042;
assign w3147 = ~w3145 & ~w3146;
assign w3148 = ~w3142 & ~w3147;
assign w3149 = ~w3143 & ~w3148;
assign w3150 = (w3149 & w2941) | (w3149 & w13830) | (w2941 & w13830);
assign w3151 = (~w2937 & w2935) | (~w2937 & w14057) | (w2935 & w14057);
assign w3152 = ~w2931 & w3151;
assign w3153 = w2937 & ~w2940;
assign w3154 = (~w3149 & w3153) | (~w3149 & w14058) | (w3153 & w14058);
assign w3155 = ~w3150 & ~w3154;
assign w3156 = ~w2728 & w3155;
assign w3157 = (~w2724 & w1570) | (~w2724 & w13831) | (w1570 & w13831);
assign w3158 = ~w1566 & w3157;
assign w3159 = (w2724 & w1571) | (w2724 & w13832) | (w1571 & w13832);
assign w3160 = ~w3158 & ~w3159;
assign w3161 = ~w3155 & ~w3160;
assign w3162 = ~w3156 & ~w3161;
assign w3163 = A_970 & A_971;
assign w3164 = A_970 & ~A_971;
assign w3165 = ~A_970 & A_971;
assign w3166 = ~w3164 & ~w3165;
assign w3167 = (~w3163 & w3166) | (~w3163 & w13514) | (w3166 & w13514);
assign w3168 = A_967 & A_968;
assign w3169 = A_967 & ~A_968;
assign w3170 = ~A_967 & A_968;
assign w3171 = ~w3169 & ~w3170;
assign w3172 = (~w3168 & w3171) | (~w3168 & w13515) | (w3171 & w13515);
assign w3173 = w3167 & ~w3172;
assign w3174 = ~w3167 & w3172;
assign w3175 = A_969 & ~w3169;
assign w3176 = ~w3170 & w3175;
assign w3177 = ~A_969 & ~w3171;
assign w3178 = ~w3176 & ~w3177;
assign w3179 = A_972 & ~w3164;
assign w3180 = ~w3165 & w3179;
assign w3181 = ~A_972 & ~w3166;
assign w3182 = ~w3180 & ~w3181;
assign w3183 = ~w3178 & ~w3182;
assign w3184 = w3183 & w3185;
assign w3185 = ~w3173 & ~w3174;
assign w3186 = ~w3183 & ~w3185;
assign w3187 = ~w3184 & ~w3186;
assign w3188 = ~w3178 & w3182;
assign w3189 = w3178 & ~w3182;
assign w3190 = ~w3188 & ~w3189;
assign w3191 = w3183 & ~w3185;
assign w3192 = ~w3167 & ~w3172;
assign w3193 = ~w3191 & ~w3192;
assign w3194 = ~w3190 & ~w3193;
assign w3195 = ~w3187 & ~w3194;
assign w3196 = ~w3187 & ~w3193;
assign w3197 = A_976 & A_977;
assign w3198 = A_976 & ~A_977;
assign w3199 = ~A_976 & A_977;
assign w3200 = ~w3198 & ~w3199;
assign w3201 = (~w3197 & w3200) | (~w3197 & w13516) | (w3200 & w13516);
assign w3202 = A_973 & A_974;
assign w3203 = A_973 & ~A_974;
assign w3204 = ~A_973 & A_974;
assign w3205 = ~w3203 & ~w3204;
assign w3206 = (~w3202 & w3205) | (~w3202 & w13517) | (w3205 & w13517);
assign w3207 = ~w3201 & w3206;
assign w3208 = w3201 & ~w3206;
assign w3209 = ~w3207 & ~w3208;
assign w3210 = A_975 & ~w3203;
assign w3211 = ~w3204 & w3210;
assign w3212 = ~A_975 & ~w3205;
assign w3213 = ~w3211 & ~w3212;
assign w3214 = A_978 & ~w3198;
assign w3215 = ~w3199 & w3214;
assign w3216 = ~A_978 & ~w3200;
assign w3217 = ~w3215 & ~w3216;
assign w3218 = ~w3213 & ~w3217;
assign w3219 = ~w3209 & w3218;
assign w3220 = ~w3201 & ~w3206;
assign w3221 = ~w3219 & ~w3220;
assign w3222 = w3218 & w3209;
assign w3223 = ~w3209 & ~w3218;
assign w3224 = ~w3222 & ~w3223;
assign w3225 = ~w3221 & ~w3224;
assign w3226 = ~w3213 & w3217;
assign w3227 = w3213 & ~w3217;
assign w3228 = ~w3226 & ~w3227;
assign w3229 = ~w3190 & ~w3228;
assign w3230 = ~w3225 & w3229;
assign w3231 = ~w3196 & w3230;
assign w3232 = ~w3221 & ~w3228;
assign w3233 = ~w3224 & ~w3232;
assign w3234 = ~w3231 & w3233;
assign w3235 = w3231 & ~w3233;
assign w3236 = ~w3234 & ~w3235;
assign w3237 = ~w3195 & ~w3236;
assign w3238 = ~w3231 & ~w3233;
assign w3239 = ~w3224 & w3229;
assign w3240 = ~w3225 & w3239;
assign w3241 = ~w3196 & ~w3232;
assign w3242 = w3240 & w3241;
assign w3243 = (w3195 & w3238) | (w3195 & w13724) | (w3238 & w13724);
assign w3244 = ~w3237 & ~w3243;
assign w3245 = A_982 & A_983;
assign w3246 = A_982 & ~A_983;
assign w3247 = ~A_982 & A_983;
assign w3248 = ~w3246 & ~w3247;
assign w3249 = (~w3245 & w3248) | (~w3245 & w13518) | (w3248 & w13518);
assign w3250 = A_979 & A_980;
assign w3251 = A_979 & ~A_980;
assign w3252 = ~A_979 & A_980;
assign w3253 = ~w3251 & ~w3252;
assign w3254 = (~w3250 & w3253) | (~w3250 & w13519) | (w3253 & w13519);
assign w3255 = w3249 & ~w3254;
assign w3256 = ~w3249 & w3254;
assign w3257 = A_981 & ~w3251;
assign w3258 = ~w3252 & w3257;
assign w3259 = ~A_981 & ~w3253;
assign w3260 = ~w3258 & ~w3259;
assign w3261 = A_984 & ~w3246;
assign w3262 = ~w3247 & w3261;
assign w3263 = ~A_984 & ~w3248;
assign w3264 = ~w3262 & ~w3263;
assign w3265 = ~w3260 & ~w3264;
assign w3266 = w3265 & w3267;
assign w3267 = ~w3255 & ~w3256;
assign w3268 = ~w3265 & ~w3267;
assign w3269 = ~w3266 & ~w3268;
assign w3270 = ~w3260 & w3264;
assign w3271 = w3260 & ~w3264;
assign w3272 = ~w3270 & ~w3271;
assign w3273 = w3265 & ~w3267;
assign w3274 = ~w3249 & ~w3254;
assign w3275 = ~w3273 & ~w3274;
assign w3276 = ~w3272 & ~w3275;
assign w3277 = ~w3269 & ~w3276;
assign w3278 = ~w3269 & ~w3275;
assign w3279 = A_988 & A_989;
assign w3280 = A_988 & ~A_989;
assign w3281 = ~A_988 & A_989;
assign w3282 = ~w3280 & ~w3281;
assign w3283 = (~w3279 & w3282) | (~w3279 & w13311) | (w3282 & w13311);
assign w3284 = A_985 & A_986;
assign w3285 = A_985 & ~A_986;
assign w3286 = ~A_985 & A_986;
assign w3287 = ~w3285 & ~w3286;
assign w3288 = (~w3284 & w3287) | (~w3284 & w13312) | (w3287 & w13312);
assign w3289 = ~w3283 & w3288;
assign w3290 = w3283 & ~w3288;
assign w3291 = ~w3289 & ~w3290;
assign w3292 = A_987 & ~w3285;
assign w3293 = ~w3286 & w3292;
assign w3294 = ~A_987 & ~w3287;
assign w3295 = ~w3293 & ~w3294;
assign w3296 = A_990 & ~w3280;
assign w3297 = ~w3281 & w3296;
assign w3298 = ~A_990 & ~w3282;
assign w3299 = ~w3297 & ~w3298;
assign w3300 = ~w3295 & ~w3299;
assign w3301 = ~w3291 & w3300;
assign w3302 = ~w3283 & ~w3288;
assign w3303 = ~w3301 & ~w3302;
assign w3304 = w3300 & w3291;
assign w3305 = ~w3291 & ~w3300;
assign w3306 = ~w3304 & ~w3305;
assign w3307 = ~w3303 & ~w3306;
assign w3308 = ~w3295 & w3299;
assign w3309 = w3295 & ~w3299;
assign w3310 = ~w3308 & ~w3309;
assign w3311 = ~w3272 & ~w3310;
assign w3312 = ~w3307 & w3311;
assign w3313 = ~w3278 & w3312;
assign w3314 = ~w3303 & ~w3310;
assign w3315 = ~w3306 & ~w3314;
assign w3316 = ~w3313 & ~w3315;
assign w3317 = ~w3306 & w3311;
assign w3318 = ~w3307 & w3317;
assign w3319 = ~w3278 & ~w3314;
assign w3320 = w3318 & w3319;
assign w3321 = (w3277 & w3316) | (w3277 & w13520) | (w3316 & w13520);
assign w3322 = ~w3313 & w3315;
assign w3323 = w3313 & ~w3315;
assign w3324 = ~w3322 & ~w3323;
assign w3325 = ~w3277 & ~w3324;
assign w3326 = ~w3307 & ~w3310;
assign w3327 = ~w3272 & ~w3278;
assign w3328 = ~w3326 & w3327;
assign w3329 = w3326 & ~w3327;
assign w3330 = ~w3328 & ~w3329;
assign w3331 = ~w3225 & ~w3228;
assign w3332 = ~w3190 & ~w3196;
assign w3333 = ~w3331 & w3332;
assign w3334 = w3331 & ~w3332;
assign w3335 = ~w3333 & ~w3334;
assign w3336 = ~w3330 & ~w3335;
assign w3337 = ~w3325 & w13725;
assign w3338 = (w3336 & w3325) | (w3336 & w13726) | (w3325 & w13726);
assign w3339 = ~w3337 & ~w3338;
assign w3340 = ~w3244 & ~w3339;
assign w3341 = ~w3325 & w13521;
assign w3342 = (~w3336 & w3325) | (~w3336 & w13727) | (w3325 & w13727);
assign w3343 = (w3244 & w3342) | (w3244 & w13522) | (w3342 & w13522);
assign w3344 = ~w3330 & w3335;
assign w3345 = w3330 & ~w3335;
assign w3346 = ~w3344 & ~w3345;
assign w3347 = ~A_961 & A_962;
assign w3348 = A_961 & ~A_962;
assign w3349 = A_963 & ~w3348;
assign w3350 = ~w3347 & w3349;
assign w3351 = ~w3347 & ~w3348;
assign w3352 = ~A_963 & ~w3351;
assign w3353 = ~w3350 & ~w3352;
assign w3354 = ~A_964 & A_965;
assign w3355 = A_964 & ~A_965;
assign w3356 = A_966 & ~w3355;
assign w3357 = ~w3354 & w3356;
assign w3358 = ~w3354 & ~w3355;
assign w3359 = ~A_966 & ~w3358;
assign w3360 = ~w3357 & ~w3359;
assign w3361 = ~w3353 & w3360;
assign w3362 = w3353 & ~w3360;
assign w3363 = ~w3361 & ~w3362;
assign w3364 = A_964 & A_965;
assign w3365 = (~w3364 & w3358) | (~w3364 & w13313) | (w3358 & w13313);
assign w3366 = A_961 & A_962;
assign w3367 = (~w3366 & w3351) | (~w3366 & w13314) | (w3351 & w13314);
assign w3368 = ~w3365 & w3367;
assign w3369 = w3365 & ~w3367;
assign w3370 = ~w3368 & ~w3369;
assign w3371 = ~w3353 & ~w3360;
assign w3372 = ~w3370 & w3371;
assign w3373 = ~w3365 & ~w3367;
assign w3374 = ~w3372 & ~w3373;
assign w3375 = w3371 & w3370;
assign w3376 = ~w3370 & ~w3371;
assign w3377 = ~w3375 & ~w3376;
assign w3378 = ~w3374 & ~w3377;
assign w3379 = ~w3363 & ~w3378;
assign w3380 = ~A_955 & A_956;
assign w3381 = A_955 & ~A_956;
assign w3382 = A_957 & ~w3381;
assign w3383 = ~w3380 & w3382;
assign w3384 = ~w3380 & ~w3381;
assign w3385 = ~A_957 & ~w3384;
assign w3386 = ~w3383 & ~w3385;
assign w3387 = ~A_958 & A_959;
assign w3388 = A_958 & ~A_959;
assign w3389 = A_960 & ~w3388;
assign w3390 = ~w3387 & w3389;
assign w3391 = ~w3387 & ~w3388;
assign w3392 = ~A_960 & ~w3391;
assign w3393 = ~w3390 & ~w3392;
assign w3394 = ~w3386 & w3393;
assign w3395 = w3386 & ~w3393;
assign w3396 = ~w3394 & ~w3395;
assign w3397 = A_958 & A_959;
assign w3398 = (~w3397 & w3391) | (~w3397 & w13523) | (w3391 & w13523);
assign w3399 = A_955 & A_956;
assign w3400 = (~w3399 & w3384) | (~w3399 & w13524) | (w3384 & w13524);
assign w3401 = ~w3398 & w3400;
assign w3402 = w3398 & ~w3400;
assign w3403 = ~w3401 & ~w3402;
assign w3404 = ~w3386 & ~w3393;
assign w3405 = ~w3403 & w3404;
assign w3406 = ~w3398 & ~w3400;
assign w3407 = ~w3405 & ~w3406;
assign w3408 = w3404 & w3403;
assign w3409 = ~w3403 & ~w3404;
assign w3410 = ~w3408 & ~w3409;
assign w3411 = ~w3407 & ~w3410;
assign w3412 = ~w3396 & ~w3411;
assign w3413 = ~w3379 & w3412;
assign w3414 = w3379 & ~w3412;
assign w3415 = ~w3413 & ~w3414;
assign w3416 = ~A_949 & A_950;
assign w3417 = A_949 & ~A_950;
assign w3418 = A_951 & ~w3417;
assign w3419 = ~w3416 & w3418;
assign w3420 = ~w3416 & ~w3417;
assign w3421 = ~A_951 & ~w3420;
assign w3422 = ~w3419 & ~w3421;
assign w3423 = ~A_952 & A_953;
assign w3424 = A_952 & ~A_953;
assign w3425 = A_954 & ~w3424;
assign w3426 = ~w3423 & w3425;
assign w3427 = ~w3423 & ~w3424;
assign w3428 = ~A_954 & ~w3427;
assign w3429 = ~w3426 & ~w3428;
assign w3430 = ~w3422 & w3429;
assign w3431 = w3422 & ~w3429;
assign w3432 = ~w3430 & ~w3431;
assign w3433 = A_952 & A_953;
assign w3434 = (~w3433 & w3427) | (~w3433 & w13525) | (w3427 & w13525);
assign w3435 = A_949 & A_950;
assign w3436 = (~w3435 & w3420) | (~w3435 & w13526) | (w3420 & w13526);
assign w3437 = ~w3434 & w3436;
assign w3438 = w3434 & ~w3436;
assign w3439 = ~w3437 & ~w3438;
assign w3440 = ~w3422 & ~w3429;
assign w3441 = ~w3439 & w3440;
assign w3442 = ~w3434 & ~w3436;
assign w3443 = ~w3441 & ~w3442;
assign w3444 = w3440 & w3439;
assign w3445 = ~w3439 & ~w3440;
assign w3446 = ~w3444 & ~w3445;
assign w3447 = ~w3443 & ~w3446;
assign w3448 = ~w3432 & ~w3447;
assign w3449 = ~A_943 & A_944;
assign w3450 = A_943 & ~A_944;
assign w3451 = A_945 & ~w3450;
assign w3452 = ~w3449 & w3451;
assign w3453 = ~w3449 & ~w3450;
assign w3454 = ~A_945 & ~w3453;
assign w3455 = ~w3452 & ~w3454;
assign w3456 = ~A_946 & A_947;
assign w3457 = A_946 & ~A_947;
assign w3458 = A_948 & ~w3457;
assign w3459 = ~w3456 & w3458;
assign w3460 = ~w3456 & ~w3457;
assign w3461 = ~A_948 & ~w3460;
assign w3462 = ~w3459 & ~w3461;
assign w3463 = ~w3455 & w3462;
assign w3464 = w3455 & ~w3462;
assign w3465 = ~w3463 & ~w3464;
assign w3466 = A_946 & A_947;
assign w3467 = (~w3466 & w3460) | (~w3466 & w13527) | (w3460 & w13527);
assign w3468 = A_943 & A_944;
assign w3469 = (~w3468 & w3453) | (~w3468 & w13528) | (w3453 & w13528);
assign w3470 = ~w3467 & w3469;
assign w3471 = w3467 & ~w3469;
assign w3472 = ~w3470 & ~w3471;
assign w3473 = ~w3455 & ~w3462;
assign w3474 = ~w3472 & w3473;
assign w3475 = ~w3467 & ~w3469;
assign w3476 = ~w3474 & ~w3475;
assign w3477 = w3473 & w3472;
assign w3478 = ~w3472 & ~w3473;
assign w3479 = ~w3477 & ~w3478;
assign w3480 = ~w3476 & ~w3479;
assign w3481 = ~w3465 & ~w3480;
assign w3482 = ~w3448 & w3481;
assign w3483 = w3448 & ~w3481;
assign w3484 = ~w3482 & ~w3483;
assign w3485 = ~w3415 & w3484;
assign w3486 = w3415 & ~w3484;
assign w3487 = ~w3485 & ~w3486;
assign w3488 = ~w3346 & ~w3487;
assign w3489 = w3488 & ~w3343;
assign w3490 = ~w3340 & w3489;
assign w3491 = ~w3340 & ~w3343;
assign w3492 = ~w3488 & ~w3491;
assign w3493 = ~w3396 & ~w3407;
assign w3494 = ~w3410 & ~w3493;
assign w3495 = ~w3363 & ~w3396;
assign w3496 = ~w3378 & w3495;
assign w3497 = ~w3411 & w3496;
assign w3498 = ~w3363 & ~w3374;
assign w3499 = ~w3377 & ~w3498;
assign w3500 = ~w3497 & ~w3499;
assign w3501 = ~w3377 & w3495;
assign w3502 = ~w3378 & w3501;
assign w3503 = ~w3411 & ~w3498;
assign w3504 = w3502 & w3503;
assign w3505 = (w3494 & w3500) | (w3494 & w13728) | (w3500 & w13728);
assign w3506 = ~w3497 & w3499;
assign w3507 = w3497 & ~w3499;
assign w3508 = ~w3506 & ~w3507;
assign w3509 = ~w3494 & ~w3508;
assign w3510 = ~w3415 & ~w3484;
assign w3511 = ~w3509 & w13729;
assign w3512 = (~w3510 & w3509) | (~w3510 & w13730) | (w3509 & w13730);
assign w3513 = ~w3511 & ~w3512;
assign w3514 = ~w3465 & ~w3476;
assign w3515 = ~w3479 & ~w3514;
assign w3516 = ~w3432 & ~w3465;
assign w3517 = ~w3447 & w3516;
assign w3518 = ~w3480 & w3517;
assign w3519 = ~w3432 & ~w3443;
assign w3520 = ~w3446 & ~w3519;
assign w3521 = ~w3518 & w3520;
assign w3522 = w3518 & ~w3520;
assign w3523 = ~w3521 & ~w3522;
assign w3524 = ~w3515 & ~w3523;
assign w3525 = ~w3518 & ~w3520;
assign w3526 = ~w3446 & w3516;
assign w3527 = ~w3447 & w3526;
assign w3528 = ~w3480 & ~w3519;
assign w3529 = w3527 & w3528;
assign w3530 = (w3515 & w3525) | (w3515 & w13833) | (w3525 & w13833);
assign w3531 = ~w3524 & ~w3530;
assign w3532 = ~w3513 & w3531;
assign w3533 = ~w3509 & w13731;
assign w3534 = (w3510 & w3509) | (w3510 & w13834) | (w3509 & w13834);
assign w3535 = (~w3531 & w3534) | (~w3531 & w13732) | (w3534 & w13732);
assign w3536 = ~w3532 & ~w3535;
assign w3537 = (w3536 & w3492) | (w3536 & w13835) | (w3492 & w13835);
assign w3538 = ~w3488 & ~w3343;
assign w3539 = ~w3340 & w3538;
assign w3540 = w3488 & ~w3491;
assign w3541 = (~w3536 & w3540) | (~w3536 & w13836) | (w3540 & w13836);
assign w3542 = ~w3537 & ~w3541;
assign w3543 = A_10 & A_11;
assign w3544 = A_10 & ~A_11;
assign w3545 = ~A_10 & A_11;
assign w3546 = ~w3544 & ~w3545;
assign w3547 = (~w3543 & w3546) | (~w3543 & w12967) | (w3546 & w12967);
assign w3548 = A_7 & A_8;
assign w3549 = A_7 & ~A_8;
assign w3550 = ~A_7 & A_8;
assign w3551 = ~w3549 & ~w3550;
assign w3552 = (~w3548 & w3551) | (~w3548 & w12968) | (w3551 & w12968);
assign w3553 = w3547 & ~w3552;
assign w3554 = ~w3547 & w3552;
assign w3555 = A_9 & ~w3549;
assign w3556 = ~w3550 & w3555;
assign w3557 = ~A_9 & ~w3551;
assign w3558 = ~w3556 & ~w3557;
assign w3559 = A_12 & ~w3544;
assign w3560 = ~w3545 & w3559;
assign w3561 = ~A_12 & ~w3546;
assign w3562 = ~w3560 & ~w3561;
assign w3563 = ~w3558 & ~w3562;
assign w3564 = w3563 & w3565;
assign w3565 = ~w3553 & ~w3554;
assign w3566 = ~w3563 & ~w3565;
assign w3567 = ~w3564 & ~w3566;
assign w3568 = ~w3558 & w3562;
assign w3569 = w3558 & ~w3562;
assign w3570 = ~w3568 & ~w3569;
assign w3571 = w3563 & ~w3565;
assign w3572 = ~w3547 & ~w3552;
assign w3573 = ~w3571 & ~w3572;
assign w3574 = ~w3570 & ~w3573;
assign w3575 = ~w3567 & ~w3574;
assign w3576 = ~w3567 & ~w3573;
assign w3577 = A_16 & A_17;
assign w3578 = A_16 & ~A_17;
assign w3579 = ~A_16 & A_17;
assign w3580 = ~w3578 & ~w3579;
assign w3581 = (~w3577 & w3580) | (~w3577 & w12704) | (w3580 & w12704);
assign w3582 = A_13 & A_14;
assign w3583 = A_13 & ~A_14;
assign w3584 = ~A_13 & A_14;
assign w3585 = ~w3583 & ~w3584;
assign w3586 = (~w3582 & w3585) | (~w3582 & w12705) | (w3585 & w12705);
assign w3587 = ~w3581 & w3586;
assign w3588 = w3581 & ~w3586;
assign w3589 = ~w3587 & ~w3588;
assign w3590 = A_15 & ~w3583;
assign w3591 = ~w3584 & w3590;
assign w3592 = ~A_15 & ~w3585;
assign w3593 = ~w3591 & ~w3592;
assign w3594 = A_18 & ~w3578;
assign w3595 = ~w3579 & w3594;
assign w3596 = ~A_18 & ~w3580;
assign w3597 = ~w3595 & ~w3596;
assign w3598 = ~w3593 & ~w3597;
assign w3599 = ~w3589 & w3598;
assign w3600 = ~w3581 & ~w3586;
assign w3601 = ~w3599 & ~w3600;
assign w3602 = w3598 & w3589;
assign w3603 = ~w3589 & ~w3598;
assign w3604 = ~w3602 & ~w3603;
assign w3605 = ~w3601 & ~w3604;
assign w3606 = ~w3593 & w3597;
assign w3607 = w3593 & ~w3597;
assign w3608 = ~w3606 & ~w3607;
assign w3609 = ~w3570 & ~w3608;
assign w3610 = ~w3605 & w3609;
assign w3611 = ~w3576 & w3610;
assign w3612 = ~w3601 & ~w3608;
assign w3613 = ~w3604 & ~w3612;
assign w3614 = ~w3611 & w3613;
assign w3615 = w3611 & ~w3613;
assign w3616 = ~w3614 & ~w3615;
assign w3617 = ~w3575 & ~w3616;
assign w3618 = ~w3611 & ~w3613;
assign w3619 = ~w3604 & w3609;
assign w3620 = ~w3605 & w3619;
assign w3621 = ~w3576 & ~w3612;
assign w3622 = w3620 & w3621;
assign w3623 = (w3575 & w3618) | (w3575 & w13315) | (w3618 & w13315);
assign w3624 = ~w3617 & ~w3623;
assign w3625 = A_22 & A_23;
assign w3626 = A_22 & ~A_23;
assign w3627 = ~A_22 & A_23;
assign w3628 = ~w3626 & ~w3627;
assign w3629 = (~w3625 & w3628) | (~w3625 & w12969) | (w3628 & w12969);
assign w3630 = A_19 & A_20;
assign w3631 = A_19 & ~A_20;
assign w3632 = ~A_19 & A_20;
assign w3633 = ~w3631 & ~w3632;
assign w3634 = (~w3630 & w3633) | (~w3630 & w12970) | (w3633 & w12970);
assign w3635 = w3629 & ~w3634;
assign w3636 = ~w3629 & w3634;
assign w3637 = A_21 & ~w3631;
assign w3638 = ~w3632 & w3637;
assign w3639 = ~A_21 & ~w3633;
assign w3640 = ~w3638 & ~w3639;
assign w3641 = A_24 & ~w3626;
assign w3642 = ~w3627 & w3641;
assign w3643 = ~A_24 & ~w3628;
assign w3644 = ~w3642 & ~w3643;
assign w3645 = ~w3640 & ~w3644;
assign w3646 = w3645 & w3647;
assign w3647 = ~w3635 & ~w3636;
assign w3648 = ~w3645 & ~w3647;
assign w3649 = ~w3646 & ~w3648;
assign w3650 = ~w3640 & w3644;
assign w3651 = w3640 & ~w3644;
assign w3652 = ~w3650 & ~w3651;
assign w3653 = w3645 & ~w3647;
assign w3654 = ~w3629 & ~w3634;
assign w3655 = ~w3653 & ~w3654;
assign w3656 = ~w3652 & ~w3655;
assign w3657 = ~w3649 & ~w3656;
assign w3658 = ~w3649 & ~w3655;
assign w3659 = A_28 & A_29;
assign w3660 = A_28 & ~A_29;
assign w3661 = ~A_28 & A_29;
assign w3662 = ~w3660 & ~w3661;
assign w3663 = (~w3659 & w3662) | (~w3659 & w12706) | (w3662 & w12706);
assign w3664 = A_25 & A_26;
assign w3665 = A_25 & ~A_26;
assign w3666 = ~A_25 & A_26;
assign w3667 = ~w3665 & ~w3666;
assign w3668 = (~w3664 & w3667) | (~w3664 & w12707) | (w3667 & w12707);
assign w3669 = ~w3663 & w3668;
assign w3670 = w3663 & ~w3668;
assign w3671 = ~w3669 & ~w3670;
assign w3672 = A_27 & ~w3665;
assign w3673 = ~w3666 & w3672;
assign w3674 = ~A_27 & ~w3667;
assign w3675 = ~w3673 & ~w3674;
assign w3676 = A_30 & ~w3660;
assign w3677 = ~w3661 & w3676;
assign w3678 = ~A_30 & ~w3662;
assign w3679 = ~w3677 & ~w3678;
assign w3680 = ~w3675 & ~w3679;
assign w3681 = ~w3671 & w3680;
assign w3682 = ~w3663 & ~w3668;
assign w3683 = ~w3681 & ~w3682;
assign w3684 = w3680 & w3671;
assign w3685 = ~w3671 & ~w3680;
assign w3686 = ~w3684 & ~w3685;
assign w3687 = ~w3683 & ~w3686;
assign w3688 = ~w3675 & w3679;
assign w3689 = w3675 & ~w3679;
assign w3690 = ~w3688 & ~w3689;
assign w3691 = ~w3652 & ~w3690;
assign w3692 = ~w3687 & w3691;
assign w3693 = ~w3658 & w3692;
assign w3694 = ~w3683 & ~w3690;
assign w3695 = ~w3686 & ~w3694;
assign w3696 = ~w3693 & ~w3695;
assign w3697 = ~w3686 & w3691;
assign w3698 = ~w3687 & w3697;
assign w3699 = ~w3658 & ~w3694;
assign w3700 = w3698 & w3699;
assign w3701 = (w3657 & w3696) | (w3657 & w12971) | (w3696 & w12971);
assign w3702 = ~w3693 & w3695;
assign w3703 = w3693 & ~w3695;
assign w3704 = ~w3702 & ~w3703;
assign w3705 = ~w3657 & ~w3704;
assign w3706 = ~w3687 & ~w3690;
assign w3707 = ~w3652 & ~w3658;
assign w3708 = ~w3706 & w3707;
assign w3709 = w3706 & ~w3707;
assign w3710 = ~w3708 & ~w3709;
assign w3711 = ~w3605 & ~w3608;
assign w3712 = ~w3570 & ~w3576;
assign w3713 = ~w3711 & w3712;
assign w3714 = w3711 & ~w3712;
assign w3715 = ~w3713 & ~w3714;
assign w3716 = ~w3710 & ~w3715;
assign w3717 = ~w3705 & w12972;
assign w3718 = (w3716 & w3705) | (w3716 & w13316) | (w3705 & w13316);
assign w3719 = ~w3717 & ~w3718;
assign w3720 = ~w3624 & ~w3719;
assign w3721 = ~w3705 & w12973;
assign w3722 = (~w3716 & w3705) | (~w3716 & w13317) | (w3705 & w13317);
assign w3723 = (w3624 & w3722) | (w3624 & w12974) | (w3722 & w12974);
assign w3724 = ~w3710 & w3715;
assign w3725 = w3710 & ~w3715;
assign w3726 = ~w3724 & ~w3725;
assign w3727 = ~A_991 & A_992;
assign w3728 = A_991 & ~A_992;
assign w3729 = A_993 & ~w3728;
assign w3730 = ~w3727 & w3729;
assign w3731 = ~w3727 & ~w3728;
assign w3732 = ~A_993 & ~w3731;
assign w3733 = ~w3730 & ~w3732;
assign w3734 = ~A_994 & A_995;
assign w3735 = A_994 & ~A_995;
assign w3736 = A_996 & ~w3735;
assign w3737 = ~w3734 & w3736;
assign w3738 = ~w3734 & ~w3735;
assign w3739 = ~A_996 & ~w3738;
assign w3740 = ~w3737 & ~w3739;
assign w3741 = ~w3733 & w3740;
assign w3742 = w3733 & ~w3740;
assign w3743 = ~w3741 & ~w3742;
assign w3744 = A_994 & A_995;
assign w3745 = (~w3744 & w3738) | (~w3744 & w13837) | (w3738 & w13837);
assign w3746 = A_991 & A_992;
assign w3747 = (~w3746 & w3731) | (~w3746 & w13838) | (w3731 & w13838);
assign w3748 = ~w3745 & w3747;
assign w3749 = w3745 & ~w3747;
assign w3750 = ~w3748 & ~w3749;
assign w3751 = ~w3733 & ~w3740;
assign w3752 = ~w3750 & w3751;
assign w3753 = ~w3745 & ~w3747;
assign w3754 = ~w3752 & ~w3753;
assign w3755 = w3751 & w3750;
assign w3756 = ~w3750 & ~w3751;
assign w3757 = ~w3755 & ~w3756;
assign w3758 = ~w3754 & ~w3757;
assign w3759 = ~w3743 & ~w3758;
assign w3760 = A_3 & ~A_4;
assign w3761 = ~A_3 & A_4;
assign w3762 = A_5 & ~w3761;
assign w3763 = ~w3760 & w3762;
assign w3764 = ~w3760 & ~w3761;
assign w3765 = ~A_5 & ~w3764;
assign w3766 = ~w3763 & ~w3765;
assign w3767 = ~A_0 & A_1;
assign w3768 = A_0 & ~A_1;
assign w3769 = ~w3767 & ~w3768;
assign w3770 = ~A_2 & ~w3769;
assign w3771 = A_2 & ~w3767;
assign w3772 = ~w3768 & w3771;
assign w3773 = (A_6 & ~w3771) | (A_6 & w12975) | (~w3771 & w12975);
assign w3774 = ~w3770 & w3773;
assign w3775 = ~w3770 & ~w3772;
assign w3776 = ~A_6 & ~w3775;
assign w3777 = (w3766 & w3776) | (w3766 & w13318) | (w3776 & w13318);
assign w3778 = ~w3766 & ~w3774;
assign w3779 = ~w3776 & w3778;
assign w3780 = ~A_997 & A_998;
assign w3781 = A_997 & ~A_998;
assign w3782 = A_999 & ~w3781;
assign w3783 = ~w3780 & w3782;
assign w3784 = ~w3780 & ~w3781;
assign w3785 = ~A_999 & ~w3784;
assign w3786 = ~w3783 & ~w3785;
assign w3787 = ~w3779 & ~w3786;
assign w3788 = ~w3777 & w3787;
assign w3789 = ~w3777 & ~w3779;
assign w3790 = w3786 & ~w3789;
assign w3791 = ~w3788 & ~w3790;
assign w3792 = w3759 & w3791;
assign w3793 = ~w3759 & ~w3791;
assign w3794 = ~w3792 & ~w3793;
assign w3795 = ~w3726 & ~w3794;
assign w3796 = w3795 & ~w3723;
assign w3797 = ~w3720 & w3796;
assign w3798 = ~w3720 & ~w3723;
assign w3799 = ~w3795 & ~w3798;
assign w3800 = ~w3743 & ~w3754;
assign w3801 = ~w3757 & ~w3800;
assign w3802 = (~w3766 & w3776) | (~w3766 & w12976) | (w3776 & w12976);
assign w3803 = A_6 & ~w3775;
assign w3804 = A_3 & A_4;
assign w3805 = (~w3804 & w3764) | (~w3804 & w13319) | (w3764 & w13319);
assign w3806 = A_0 & A_1;
assign w3807 = (~w3806 & w3769) | (~w3806 & w13320) | (w3769 & w13320);
assign w3808 = ~w3805 & w3807;
assign w3809 = w3805 & ~w3807;
assign w3810 = ~w3808 & ~w3809;
assign w3811 = ~w3803 & w3810;
assign w3812 = ~w3802 & w3811;
assign w3813 = (~w3810 & w3802) | (~w3810 & w13321) | (w3802 & w13321);
assign w3814 = ~w3812 & ~w3813;
assign w3815 = ~w3786 & ~w3789;
assign w3816 = w3814 & w3815;
assign w3817 = A_997 & A_998;
assign w3818 = (~w3817 & w3784) | (~w3817 & w13839) | (w3784 & w13839);
assign w3819 = ~w3814 & ~w3815;
assign w3820 = w3818 & ~w3819;
assign w3821 = ~w3816 & w3820;
assign w3822 = ~w3816 & ~w3819;
assign w3823 = ~w3818 & ~w3822;
assign w3824 = w3759 & ~w3791;
assign w3825 = ~w3823 & w3824;
assign w3826 = ~w3821 & w3825;
assign w3827 = ~w3821 & ~w3823;
assign w3828 = ~w3824 & ~w3827;
assign w3829 = ~w3826 & ~w3828;
assign w3830 = ~w3801 & ~w3829;
assign w3831 = ~w3823 & ~w3824;
assign w3832 = ~w3821 & w3831;
assign w3833 = w3824 & ~w3827;
assign w3834 = ~w3832 & ~w3833;
assign w3835 = w3801 & ~w3834;
assign w3836 = ~w3830 & ~w3835;
assign w3837 = (w3836 & w3799) | (w3836 & w13840) | (w3799 & w13840);
assign w3838 = ~w3795 & ~w3723;
assign w3839 = ~w3720 & w3838;
assign w3840 = w3795 & ~w3798;
assign w3841 = (~w3836 & w3840) | (~w3836 & w13841) | (w3840 & w13841);
assign w3842 = ~w3837 & ~w3841;
assign w3843 = A_46 & A_47;
assign w3844 = A_46 & ~A_47;
assign w3845 = ~A_46 & A_47;
assign w3846 = ~w3844 & ~w3845;
assign w3847 = (~w3843 & w3846) | (~w3843 & w12708) | (w3846 & w12708);
assign w3848 = A_43 & A_44;
assign w3849 = A_43 & ~A_44;
assign w3850 = ~A_43 & A_44;
assign w3851 = ~w3849 & ~w3850;
assign w3852 = (~w3848 & w3851) | (~w3848 & w12709) | (w3851 & w12709);
assign w3853 = w3847 & ~w3852;
assign w3854 = ~w3847 & w3852;
assign w3855 = A_45 & ~w3849;
assign w3856 = ~w3850 & w3855;
assign w3857 = ~A_45 & ~w3851;
assign w3858 = ~w3856 & ~w3857;
assign w3859 = A_48 & ~w3844;
assign w3860 = ~w3845 & w3859;
assign w3861 = ~A_48 & ~w3846;
assign w3862 = ~w3860 & ~w3861;
assign w3863 = ~w3858 & ~w3862;
assign w3864 = w3863 & w3865;
assign w3865 = ~w3853 & ~w3854;
assign w3866 = ~w3863 & ~w3865;
assign w3867 = ~w3864 & ~w3866;
assign w3868 = ~w3858 & w3862;
assign w3869 = w3858 & ~w3862;
assign w3870 = ~w3868 & ~w3869;
assign w3871 = w3863 & ~w3865;
assign w3872 = ~w3847 & ~w3852;
assign w3873 = ~w3871 & ~w3872;
assign w3874 = ~w3870 & ~w3873;
assign w3875 = ~w3867 & ~w3874;
assign w3876 = ~w3867 & ~w3873;
assign w3877 = A_52 & A_53;
assign w3878 = A_52 & ~A_53;
assign w3879 = ~A_52 & A_53;
assign w3880 = ~w3878 & ~w3879;
assign w3881 = (~w3877 & w3880) | (~w3877 & w12710) | (w3880 & w12710);
assign w3882 = A_49 & A_50;
assign w3883 = A_49 & ~A_50;
assign w3884 = ~A_49 & A_50;
assign w3885 = ~w3883 & ~w3884;
assign w3886 = (~w3882 & w3885) | (~w3882 & w12711) | (w3885 & w12711);
assign w3887 = ~w3881 & w3886;
assign w3888 = w3881 & ~w3886;
assign w3889 = ~w3887 & ~w3888;
assign w3890 = A_51 & ~w3883;
assign w3891 = ~w3884 & w3890;
assign w3892 = ~A_51 & ~w3885;
assign w3893 = ~w3891 & ~w3892;
assign w3894 = A_54 & ~w3878;
assign w3895 = ~w3879 & w3894;
assign w3896 = ~A_54 & ~w3880;
assign w3897 = ~w3895 & ~w3896;
assign w3898 = ~w3893 & ~w3897;
assign w3899 = ~w3889 & w3898;
assign w3900 = ~w3881 & ~w3886;
assign w3901 = ~w3899 & ~w3900;
assign w3902 = w3898 & w3889;
assign w3903 = ~w3889 & ~w3898;
assign w3904 = ~w3902 & ~w3903;
assign w3905 = ~w3901 & ~w3904;
assign w3906 = ~w3893 & w3897;
assign w3907 = w3893 & ~w3897;
assign w3908 = ~w3906 & ~w3907;
assign w3909 = ~w3870 & ~w3908;
assign w3910 = ~w3905 & w3909;
assign w3911 = ~w3876 & w3910;
assign w3912 = ~w3901 & ~w3908;
assign w3913 = ~w3904 & ~w3912;
assign w3914 = ~w3911 & ~w3913;
assign w3915 = ~w3904 & w3909;
assign w3916 = ~w3905 & w3915;
assign w3917 = ~w3876 & ~w3912;
assign w3918 = w3916 & w3917;
assign w3919 = (w3875 & w3914) | (w3875 & w12977) | (w3914 & w12977);
assign w3920 = ~w3911 & w3913;
assign w3921 = w3911 & ~w3913;
assign w3922 = ~w3920 & ~w3921;
assign w3923 = ~w3875 & ~w3922;
assign w3924 = ~w3905 & ~w3908;
assign w3925 = ~w3870 & ~w3876;
assign w3926 = ~w3924 & w3925;
assign w3927 = w3924 & ~w3925;
assign w3928 = ~w3926 & ~w3927;
assign w3929 = ~A_37 & A_38;
assign w3930 = A_37 & ~A_38;
assign w3931 = A_39 & ~w3930;
assign w3932 = ~w3929 & w3931;
assign w3933 = ~w3929 & ~w3930;
assign w3934 = ~A_39 & ~w3933;
assign w3935 = ~w3932 & ~w3934;
assign w3936 = ~A_40 & A_41;
assign w3937 = A_40 & ~A_41;
assign w3938 = A_42 & ~w3937;
assign w3939 = ~w3936 & w3938;
assign w3940 = ~w3936 & ~w3937;
assign w3941 = ~A_42 & ~w3940;
assign w3942 = ~w3939 & ~w3941;
assign w3943 = ~w3935 & w3942;
assign w3944 = w3935 & ~w3942;
assign w3945 = ~w3943 & ~w3944;
assign w3946 = A_40 & A_41;
assign w3947 = (~w3946 & w3940) | (~w3946 & w12712) | (w3940 & w12712);
assign w3948 = A_37 & A_38;
assign w3949 = (~w3948 & w3933) | (~w3948 & w12713) | (w3933 & w12713);
assign w3950 = ~w3947 & w3949;
assign w3951 = w3947 & ~w3949;
assign w3952 = ~w3950 & ~w3951;
assign w3953 = ~w3935 & ~w3942;
assign w3954 = ~w3952 & w3953;
assign w3955 = ~w3947 & ~w3949;
assign w3956 = ~w3954 & ~w3955;
assign w3957 = w3953 & w3952;
assign w3958 = ~w3952 & ~w3953;
assign w3959 = ~w3957 & ~w3958;
assign w3960 = ~w3956 & ~w3959;
assign w3961 = ~w3945 & ~w3960;
assign w3962 = ~A_31 & A_32;
assign w3963 = A_31 & ~A_32;
assign w3964 = A_33 & ~w3963;
assign w3965 = ~w3962 & w3964;
assign w3966 = ~w3962 & ~w3963;
assign w3967 = ~A_33 & ~w3966;
assign w3968 = ~w3965 & ~w3967;
assign w3969 = ~A_34 & A_35;
assign w3970 = A_34 & ~A_35;
assign w3971 = A_36 & ~w3970;
assign w3972 = ~w3969 & w3971;
assign w3973 = ~w3969 & ~w3970;
assign w3974 = ~A_36 & ~w3973;
assign w3975 = ~w3972 & ~w3974;
assign w3976 = ~w3968 & w3975;
assign w3977 = w3968 & ~w3975;
assign w3978 = ~w3976 & ~w3977;
assign w3979 = A_34 & A_35;
assign w3980 = (~w3979 & w3973) | (~w3979 & w12714) | (w3973 & w12714);
assign w3981 = A_31 & A_32;
assign w3982 = (~w3981 & w3966) | (~w3981 & w12715) | (w3966 & w12715);
assign w3983 = ~w3980 & w3982;
assign w3984 = w3980 & ~w3982;
assign w3985 = ~w3983 & ~w3984;
assign w3986 = ~w3968 & ~w3975;
assign w3987 = ~w3985 & w3986;
assign w3988 = ~w3980 & ~w3982;
assign w3989 = ~w3987 & ~w3988;
assign w3990 = w3986 & w3985;
assign w3991 = ~w3985 & ~w3986;
assign w3992 = ~w3990 & ~w3991;
assign w3993 = ~w3989 & ~w3992;
assign w3994 = ~w3978 & ~w3993;
assign w3995 = ~w3961 & w3994;
assign w3996 = w3961 & ~w3994;
assign w3997 = ~w3995 & ~w3996;
assign w3998 = ~w3928 & ~w3997;
assign w3999 = ~w3923 & w13322;
assign w4000 = (~w3998 & w3923) | (~w3998 & w13323) | (w3923 & w13323);
assign w4001 = ~w3999 & ~w4000;
assign w4002 = ~w3978 & ~w3989;
assign w4003 = ~w3992 & ~w4002;
assign w4004 = ~w3945 & ~w3978;
assign w4005 = ~w3960 & w4004;
assign w4006 = ~w3993 & w4005;
assign w4007 = ~w3945 & ~w3956;
assign w4008 = ~w3959 & ~w4007;
assign w4009 = ~w4006 & w4008;
assign w4010 = w4006 & ~w4008;
assign w4011 = ~w4009 & ~w4010;
assign w4012 = ~w4003 & ~w4011;
assign w4013 = ~w4006 & ~w4008;
assign w4014 = ~w3959 & w4004;
assign w4015 = ~w3960 & w4014;
assign w4016 = ~w3993 & ~w4007;
assign w4017 = w4015 & w4016;
assign w4018 = (w4003 & w4013) | (w4003 & w13324) | (w4013 & w13324);
assign w4019 = ~w4012 & ~w4018;
assign w4020 = ~w4001 & w4019;
assign w4021 = ~w3923 & w12978;
assign w4022 = (w3998 & w3923) | (w3998 & w13325) | (w3923 & w13325);
assign w4023 = ~w4021 & ~w4022;
assign w4024 = ~w4019 & ~w4023;
assign w4025 = ~w4020 & ~w4024;
assign w4026 = A_58 & A_59;
assign w4027 = A_58 & ~A_59;
assign w4028 = ~A_58 & A_59;
assign w4029 = ~w4027 & ~w4028;
assign w4030 = (~w4026 & w4029) | (~w4026 & w12716) | (w4029 & w12716);
assign w4031 = A_55 & A_56;
assign w4032 = A_55 & ~A_56;
assign w4033 = ~A_55 & A_56;
assign w4034 = ~w4032 & ~w4033;
assign w4035 = (~w4031 & w4034) | (~w4031 & w12717) | (w4034 & w12717);
assign w4036 = w4030 & ~w4035;
assign w4037 = ~w4030 & w4035;
assign w4038 = A_57 & ~w4032;
assign w4039 = ~w4033 & w4038;
assign w4040 = ~A_57 & ~w4034;
assign w4041 = ~w4039 & ~w4040;
assign w4042 = A_60 & ~w4027;
assign w4043 = ~w4028 & w4042;
assign w4044 = ~A_60 & ~w4029;
assign w4045 = ~w4043 & ~w4044;
assign w4046 = ~w4041 & ~w4045;
assign w4047 = w4046 & w4048;
assign w4048 = ~w4036 & ~w4037;
assign w4049 = ~w4046 & ~w4048;
assign w4050 = ~w4047 & ~w4049;
assign w4051 = ~w4041 & w4045;
assign w4052 = w4041 & ~w4045;
assign w4053 = ~w4051 & ~w4052;
assign w4054 = w4046 & ~w4048;
assign w4055 = ~w4030 & ~w4035;
assign w4056 = ~w4054 & ~w4055;
assign w4057 = ~w4053 & ~w4056;
assign w4058 = ~w4050 & ~w4057;
assign w4059 = ~w4050 & ~w4056;
assign w4060 = A_64 & A_65;
assign w4061 = A_64 & ~A_65;
assign w4062 = ~A_64 & A_65;
assign w4063 = ~w4061 & ~w4062;
assign w4064 = (~w4060 & w4063) | (~w4060 & w12718) | (w4063 & w12718);
assign w4065 = A_61 & A_62;
assign w4066 = A_61 & ~A_62;
assign w4067 = ~A_61 & A_62;
assign w4068 = ~w4066 & ~w4067;
assign w4069 = (~w4065 & w4068) | (~w4065 & w12719) | (w4068 & w12719);
assign w4070 = ~w4064 & w4069;
assign w4071 = w4064 & ~w4069;
assign w4072 = ~w4070 & ~w4071;
assign w4073 = A_63 & ~w4066;
assign w4074 = ~w4067 & w4073;
assign w4075 = ~A_63 & ~w4068;
assign w4076 = ~w4074 & ~w4075;
assign w4077 = A_66 & ~w4061;
assign w4078 = ~w4062 & w4077;
assign w4079 = ~A_66 & ~w4063;
assign w4080 = ~w4078 & ~w4079;
assign w4081 = ~w4076 & ~w4080;
assign w4082 = ~w4072 & w4081;
assign w4083 = ~w4064 & ~w4069;
assign w4084 = ~w4082 & ~w4083;
assign w4085 = w4081 & w4072;
assign w4086 = ~w4072 & ~w4081;
assign w4087 = ~w4085 & ~w4086;
assign w4088 = ~w4084 & ~w4087;
assign w4089 = ~w4076 & w4080;
assign w4090 = w4076 & ~w4080;
assign w4091 = ~w4089 & ~w4090;
assign w4092 = ~w4053 & ~w4091;
assign w4093 = ~w4088 & w4092;
assign w4094 = ~w4059 & w4093;
assign w4095 = ~w4084 & ~w4091;
assign w4096 = ~w4087 & ~w4095;
assign w4097 = ~w4094 & w4096;
assign w4098 = w4094 & ~w4096;
assign w4099 = ~w4097 & ~w4098;
assign w4100 = ~w4058 & ~w4099;
assign w4101 = ~w4094 & ~w4096;
assign w4102 = ~w4087 & w4092;
assign w4103 = ~w4088 & w4102;
assign w4104 = ~w4059 & ~w4095;
assign w4105 = w4103 & w4104;
assign w4106 = (w4058 & w4101) | (w4058 & w13326) | (w4101 & w13326);
assign w4107 = ~w4100 & ~w4106;
assign w4108 = A_70 & A_71;
assign w4109 = A_70 & ~A_71;
assign w4110 = ~A_70 & A_71;
assign w4111 = ~w4109 & ~w4110;
assign w4112 = (~w4108 & w4111) | (~w4108 & w12720) | (w4111 & w12720);
assign w4113 = A_67 & A_68;
assign w4114 = A_67 & ~A_68;
assign w4115 = ~A_67 & A_68;
assign w4116 = ~w4114 & ~w4115;
assign w4117 = (~w4113 & w4116) | (~w4113 & w12721) | (w4116 & w12721);
assign w4118 = w4112 & ~w4117;
assign w4119 = ~w4112 & w4117;
assign w4120 = A_69 & ~w4114;
assign w4121 = ~w4115 & w4120;
assign w4122 = ~A_69 & ~w4116;
assign w4123 = ~w4121 & ~w4122;
assign w4124 = A_72 & ~w4109;
assign w4125 = ~w4110 & w4124;
assign w4126 = ~A_72 & ~w4111;
assign w4127 = ~w4125 & ~w4126;
assign w4128 = ~w4123 & ~w4127;
assign w4129 = w4128 & w4130;
assign w4130 = ~w4118 & ~w4119;
assign w4131 = ~w4128 & ~w4130;
assign w4132 = ~w4129 & ~w4131;
assign w4133 = ~w4123 & w4127;
assign w4134 = w4123 & ~w4127;
assign w4135 = ~w4133 & ~w4134;
assign w4136 = w4128 & ~w4130;
assign w4137 = ~w4112 & ~w4117;
assign w4138 = ~w4136 & ~w4137;
assign w4139 = ~w4135 & ~w4138;
assign w4140 = ~w4132 & ~w4139;
assign w4141 = ~w4132 & ~w4138;
assign w4142 = A_76 & A_77;
assign w4143 = A_76 & ~A_77;
assign w4144 = ~A_76 & A_77;
assign w4145 = ~w4143 & ~w4144;
assign w4146 = (~w4142 & w4145) | (~w4142 & w12722) | (w4145 & w12722);
assign w4147 = A_73 & A_74;
assign w4148 = A_73 & ~A_74;
assign w4149 = ~A_73 & A_74;
assign w4150 = ~w4148 & ~w4149;
assign w4151 = (~w4147 & w4150) | (~w4147 & w12723) | (w4150 & w12723);
assign w4152 = ~w4146 & w4151;
assign w4153 = w4146 & ~w4151;
assign w4154 = ~w4152 & ~w4153;
assign w4155 = A_75 & ~w4148;
assign w4156 = ~w4149 & w4155;
assign w4157 = ~A_75 & ~w4150;
assign w4158 = ~w4156 & ~w4157;
assign w4159 = A_78 & ~w4143;
assign w4160 = ~w4144 & w4159;
assign w4161 = ~A_78 & ~w4145;
assign w4162 = ~w4160 & ~w4161;
assign w4163 = ~w4158 & ~w4162;
assign w4164 = ~w4154 & w4163;
assign w4165 = ~w4146 & ~w4151;
assign w4166 = ~w4164 & ~w4165;
assign w4167 = w4163 & w4154;
assign w4168 = ~w4154 & ~w4163;
assign w4169 = ~w4167 & ~w4168;
assign w4170 = ~w4166 & ~w4169;
assign w4171 = ~w4158 & w4162;
assign w4172 = w4158 & ~w4162;
assign w4173 = ~w4171 & ~w4172;
assign w4174 = ~w4135 & ~w4173;
assign w4175 = ~w4170 & w4174;
assign w4176 = ~w4141 & w4175;
assign w4177 = ~w4166 & ~w4173;
assign w4178 = ~w4169 & ~w4177;
assign w4179 = ~w4176 & ~w4178;
assign w4180 = ~w4169 & w4174;
assign w4181 = ~w4170 & w4180;
assign w4182 = ~w4141 & ~w4177;
assign w4183 = w4181 & w4182;
assign w4184 = (w4140 & w4179) | (w4140 & w12979) | (w4179 & w12979);
assign w4185 = ~w4176 & w4178;
assign w4186 = w4176 & ~w4178;
assign w4187 = ~w4185 & ~w4186;
assign w4188 = ~w4140 & ~w4187;
assign w4189 = ~w4170 & ~w4173;
assign w4190 = ~w4135 & ~w4141;
assign w4191 = ~w4189 & w4190;
assign w4192 = w4189 & ~w4190;
assign w4193 = ~w4191 & ~w4192;
assign w4194 = ~w4088 & ~w4091;
assign w4195 = ~w4053 & ~w4059;
assign w4196 = ~w4194 & w4195;
assign w4197 = w4194 & ~w4195;
assign w4198 = ~w4196 & ~w4197;
assign w4199 = ~w4193 & ~w4198;
assign w4200 = ~w4188 & w12980;
assign w4201 = (w4199 & w4188) | (w4199 & w12981) | (w4188 & w12981);
assign w4202 = ~w4200 & ~w4201;
assign w4203 = ~w4107 & ~w4202;
assign w4204 = ~w4188 & w12982;
assign w4205 = (~w4199 & w4188) | (~w4199 & w13327) | (w4188 & w13327);
assign w4206 = (w4107 & w4205) | (w4107 & w12983) | (w4205 & w12983);
assign w4207 = ~w4193 & w4198;
assign w4208 = w4193 & ~w4198;
assign w4209 = ~w4207 & ~w4208;
assign w4210 = ~w3928 & w3997;
assign w4211 = w3928 & ~w3997;
assign w4212 = ~w4210 & ~w4211;
assign w4213 = ~w4209 & ~w4212;
assign w4214 = ~w4213 & ~w4206;
assign w4215 = ~w4203 & w4214;
assign w4216 = ~w4203 & ~w4206;
assign w4217 = w4213 & ~w4216;
assign w4218 = (~w4025 & w4217) | (~w4025 & w13328) | (w4217 & w13328);
assign w4219 = w4213 & ~w4206;
assign w4220 = ~w4203 & w4219;
assign w4221 = ~w4213 & ~w4216;
assign w4222 = ~w4220 & ~w4221;
assign w4223 = (w4025 & w4221) | (w4025 & w13842) | (w4221 & w13842);
assign w4224 = ~w4209 & w4212;
assign w4225 = w4209 & ~w4212;
assign w4226 = ~w4224 & ~w4225;
assign w4227 = ~w3726 & w3794;
assign w4228 = ~w3724 & ~w3794;
assign w4229 = ~w3725 & w4228;
assign w4230 = ~w4227 & ~w4229;
assign w4231 = ~w4226 & ~w4230;
assign w4232 = (~w4231 & w4222) | (~w4231 & w13329) | (w4222 & w13329);
assign w4233 = ~w4218 & w4232;
assign w4234 = (w4231 & w4223) | (w4231 & w13330) | (w4223 & w13330);
assign w4235 = ~w4233 & ~w4234;
assign w4236 = ~w3842 & ~w4235;
assign w4237 = (w4231 & w4222) | (w4231 & w13331) | (w4222 & w13331);
assign w4238 = ~w4218 & w4237;
assign w4239 = (~w4231 & w4223) | (~w4231 & w13332) | (w4223 & w13332);
assign w4240 = ~w4238 & ~w4239;
assign w4241 = w3842 & ~w4240;
assign w4242 = ~w4226 & w4230;
assign w4243 = w4226 & ~w4230;
assign w4244 = ~w4242 & ~w4243;
assign w4245 = ~w3346 & w3487;
assign w4246 = w3346 & ~w3487;
assign w4247 = ~w4245 & ~w4246;
assign w4248 = ~w4244 & ~w4247;
assign w4249 = (~w4248 & w4240) | (~w4248 & w13843) | (w4240 & w13843);
assign w4250 = ~w4236 & w4249;
assign w4251 = ~w4236 & ~w4241;
assign w4252 = w4248 & ~w4251;
assign w4253 = ~w4250 & ~w4252;
assign w4254 = (~w3542 & w4252) | (~w3542 & w13844) | (w4252 & w13844);
assign w4255 = (w4248 & w4240) | (w4248 & w13845) | (w4240 & w13845);
assign w4256 = ~w4236 & w4255;
assign w4257 = ~w4248 & ~w4251;
assign w4258 = (w3542 & w4257) | (w3542 & w13846) | (w4257 & w13846);
assign w4259 = ~w4244 & w4247;
assign w4260 = ~w4242 & ~w4247;
assign w4261 = ~w4243 & w4260;
assign w4262 = ~w4259 & ~w4261;
assign w4263 = ~A_937 & A_938;
assign w4264 = A_937 & ~A_938;
assign w4265 = A_939 & ~w4264;
assign w4266 = ~w4263 & w4265;
assign w4267 = ~w4263 & ~w4264;
assign w4268 = ~A_939 & ~w4267;
assign w4269 = ~w4266 & ~w4268;
assign w4270 = ~A_940 & A_941;
assign w4271 = A_940 & ~A_941;
assign w4272 = A_942 & ~w4271;
assign w4273 = ~w4270 & w4272;
assign w4274 = ~w4270 & ~w4271;
assign w4275 = ~A_942 & ~w4274;
assign w4276 = ~w4273 & ~w4275;
assign w4277 = ~w4269 & w4276;
assign w4278 = w4269 & ~w4276;
assign w4279 = ~w4277 & ~w4278;
assign w4280 = A_940 & A_941;
assign w4281 = (~w4280 & w4274) | (~w4280 & w13333) | (w4274 & w13333);
assign w4282 = A_937 & A_938;
assign w4283 = (~w4282 & w4267) | (~w4282 & w13334) | (w4267 & w13334);
assign w4284 = ~w4281 & w4283;
assign w4285 = w4281 & ~w4283;
assign w4286 = ~w4284 & ~w4285;
assign w4287 = ~w4269 & ~w4276;
assign w4288 = ~w4286 & w4287;
assign w4289 = ~w4281 & ~w4283;
assign w4290 = ~w4288 & ~w4289;
assign w4291 = w4287 & w4286;
assign w4292 = ~w4286 & ~w4287;
assign w4293 = ~w4291 & ~w4292;
assign w4294 = ~w4290 & ~w4293;
assign w4295 = ~w4279 & ~w4294;
assign w4296 = ~A_931 & A_932;
assign w4297 = A_931 & ~A_932;
assign w4298 = A_933 & ~w4297;
assign w4299 = ~w4296 & w4298;
assign w4300 = ~w4296 & ~w4297;
assign w4301 = ~A_933 & ~w4300;
assign w4302 = ~w4299 & ~w4301;
assign w4303 = ~A_934 & A_935;
assign w4304 = A_934 & ~A_935;
assign w4305 = A_936 & ~w4304;
assign w4306 = ~w4303 & w4305;
assign w4307 = ~w4303 & ~w4304;
assign w4308 = ~A_936 & ~w4307;
assign w4309 = ~w4306 & ~w4308;
assign w4310 = ~w4302 & w4309;
assign w4311 = w4302 & ~w4309;
assign w4312 = ~w4310 & ~w4311;
assign w4313 = A_934 & A_935;
assign w4314 = (~w4313 & w4307) | (~w4313 & w13335) | (w4307 & w13335);
assign w4315 = A_931 & A_932;
assign w4316 = (~w4315 & w4300) | (~w4315 & w13336) | (w4300 & w13336);
assign w4317 = ~w4314 & w4316;
assign w4318 = w4314 & ~w4316;
assign w4319 = ~w4317 & ~w4318;
assign w4320 = ~w4302 & ~w4309;
assign w4321 = ~w4319 & w4320;
assign w4322 = ~w4314 & ~w4316;
assign w4323 = ~w4321 & ~w4322;
assign w4324 = w4320 & w4319;
assign w4325 = ~w4319 & ~w4320;
assign w4326 = ~w4324 & ~w4325;
assign w4327 = ~w4323 & ~w4326;
assign w4328 = ~w4312 & ~w4327;
assign w4329 = ~w4295 & w4328;
assign w4330 = w4295 & ~w4328;
assign w4331 = ~w4329 & ~w4330;
assign w4332 = ~A_925 & A_926;
assign w4333 = A_925 & ~A_926;
assign w4334 = A_927 & ~w4333;
assign w4335 = ~w4332 & w4334;
assign w4336 = ~w4332 & ~w4333;
assign w4337 = ~A_927 & ~w4336;
assign w4338 = ~w4335 & ~w4337;
assign w4339 = ~A_928 & A_929;
assign w4340 = A_928 & ~A_929;
assign w4341 = A_930 & ~w4340;
assign w4342 = ~w4339 & w4341;
assign w4343 = ~w4339 & ~w4340;
assign w4344 = ~A_930 & ~w4343;
assign w4345 = ~w4342 & ~w4344;
assign w4346 = ~w4338 & w4345;
assign w4347 = w4338 & ~w4345;
assign w4348 = ~w4346 & ~w4347;
assign w4349 = A_928 & A_929;
assign w4350 = (~w4349 & w4343) | (~w4349 & w13337) | (w4343 & w13337);
assign w4351 = A_925 & A_926;
assign w4352 = (~w4351 & w4336) | (~w4351 & w13338) | (w4336 & w13338);
assign w4353 = ~w4350 & w4352;
assign w4354 = w4350 & ~w4352;
assign w4355 = ~w4353 & ~w4354;
assign w4356 = ~w4338 & ~w4345;
assign w4357 = ~w4355 & w4356;
assign w4358 = ~w4350 & ~w4352;
assign w4359 = ~w4357 & ~w4358;
assign w4360 = w4356 & w4355;
assign w4361 = ~w4355 & ~w4356;
assign w4362 = ~w4360 & ~w4361;
assign w4363 = ~w4359 & ~w4362;
assign w4364 = ~w4348 & ~w4363;
assign w4365 = ~A_919 & A_920;
assign w4366 = A_919 & ~A_920;
assign w4367 = A_921 & ~w4366;
assign w4368 = ~w4365 & w4367;
assign w4369 = ~w4365 & ~w4366;
assign w4370 = ~A_921 & ~w4369;
assign w4371 = ~w4368 & ~w4370;
assign w4372 = ~A_922 & A_923;
assign w4373 = A_922 & ~A_923;
assign w4374 = A_924 & ~w4373;
assign w4375 = ~w4372 & w4374;
assign w4376 = ~w4372 & ~w4373;
assign w4377 = ~A_924 & ~w4376;
assign w4378 = ~w4375 & ~w4377;
assign w4379 = ~w4371 & w4378;
assign w4380 = w4371 & ~w4378;
assign w4381 = ~w4379 & ~w4380;
assign w4382 = A_922 & A_923;
assign w4383 = (~w4382 & w4376) | (~w4382 & w13339) | (w4376 & w13339);
assign w4384 = A_919 & A_920;
assign w4385 = (~w4384 & w4369) | (~w4384 & w13340) | (w4369 & w13340);
assign w4386 = ~w4383 & w4385;
assign w4387 = w4383 & ~w4385;
assign w4388 = ~w4386 & ~w4387;
assign w4389 = ~w4371 & ~w4378;
assign w4390 = ~w4388 & w4389;
assign w4391 = ~w4383 & ~w4385;
assign w4392 = ~w4390 & ~w4391;
assign w4393 = w4389 & w4388;
assign w4394 = ~w4388 & ~w4389;
assign w4395 = ~w4393 & ~w4394;
assign w4396 = ~w4392 & ~w4395;
assign w4397 = ~w4381 & ~w4396;
assign w4398 = ~w4364 & w4397;
assign w4399 = w4364 & ~w4397;
assign w4400 = ~w4398 & ~w4399;
assign w4401 = ~w4331 & w4400;
assign w4402 = w4331 & ~w4400;
assign w4403 = ~w4401 & ~w4402;
assign w4404 = ~A_913 & A_914;
assign w4405 = A_913 & ~A_914;
assign w4406 = A_915 & ~w4405;
assign w4407 = ~w4404 & w4406;
assign w4408 = ~w4404 & ~w4405;
assign w4409 = ~A_915 & ~w4408;
assign w4410 = ~w4407 & ~w4409;
assign w4411 = ~A_916 & A_917;
assign w4412 = A_916 & ~A_917;
assign w4413 = A_918 & ~w4412;
assign w4414 = ~w4411 & w4413;
assign w4415 = ~w4411 & ~w4412;
assign w4416 = ~A_918 & ~w4415;
assign w4417 = ~w4414 & ~w4416;
assign w4418 = ~w4410 & w4417;
assign w4419 = w4410 & ~w4417;
assign w4420 = ~w4418 & ~w4419;
assign w4421 = A_916 & A_917;
assign w4422 = (~w4421 & w4415) | (~w4421 & w13341) | (w4415 & w13341);
assign w4423 = A_913 & A_914;
assign w4424 = (~w4423 & w4408) | (~w4423 & w13342) | (w4408 & w13342);
assign w4425 = ~w4422 & w4424;
assign w4426 = w4422 & ~w4424;
assign w4427 = ~w4425 & ~w4426;
assign w4428 = ~w4410 & ~w4417;
assign w4429 = ~w4427 & w4428;
assign w4430 = ~w4422 & ~w4424;
assign w4431 = ~w4429 & ~w4430;
assign w4432 = w4428 & w4427;
assign w4433 = ~w4427 & ~w4428;
assign w4434 = ~w4432 & ~w4433;
assign w4435 = ~w4431 & ~w4434;
assign w4436 = ~w4420 & ~w4435;
assign w4437 = ~A_907 & A_908;
assign w4438 = A_907 & ~A_908;
assign w4439 = A_909 & ~w4438;
assign w4440 = ~w4437 & w4439;
assign w4441 = ~w4437 & ~w4438;
assign w4442 = ~A_909 & ~w4441;
assign w4443 = ~w4440 & ~w4442;
assign w4444 = ~A_910 & A_911;
assign w4445 = A_910 & ~A_911;
assign w4446 = A_912 & ~w4445;
assign w4447 = ~w4444 & w4446;
assign w4448 = ~w4444 & ~w4445;
assign w4449 = ~A_912 & ~w4448;
assign w4450 = ~w4447 & ~w4449;
assign w4451 = ~w4443 & w4450;
assign w4452 = w4443 & ~w4450;
assign w4453 = ~w4451 & ~w4452;
assign w4454 = A_910 & A_911;
assign w4455 = (~w4454 & w4448) | (~w4454 & w13343) | (w4448 & w13343);
assign w4456 = A_907 & A_908;
assign w4457 = (~w4456 & w4441) | (~w4456 & w13344) | (w4441 & w13344);
assign w4458 = ~w4455 & w4457;
assign w4459 = w4455 & ~w4457;
assign w4460 = ~w4458 & ~w4459;
assign w4461 = ~w4443 & ~w4450;
assign w4462 = ~w4460 & w4461;
assign w4463 = ~w4455 & ~w4457;
assign w4464 = ~w4462 & ~w4463;
assign w4465 = w4461 & w4460;
assign w4466 = ~w4460 & ~w4461;
assign w4467 = ~w4465 & ~w4466;
assign w4468 = ~w4464 & ~w4467;
assign w4469 = ~w4453 & ~w4468;
assign w4470 = ~w4436 & w4469;
assign w4471 = w4436 & ~w4469;
assign w4472 = ~w4470 & ~w4471;
assign w4473 = ~A_901 & A_902;
assign w4474 = A_901 & ~A_902;
assign w4475 = A_903 & ~w4474;
assign w4476 = ~w4473 & w4475;
assign w4477 = ~w4473 & ~w4474;
assign w4478 = ~A_903 & ~w4477;
assign w4479 = ~w4476 & ~w4478;
assign w4480 = ~A_904 & A_905;
assign w4481 = A_904 & ~A_905;
assign w4482 = A_906 & ~w4481;
assign w4483 = ~w4480 & w4482;
assign w4484 = ~w4480 & ~w4481;
assign w4485 = ~A_906 & ~w4484;
assign w4486 = ~w4483 & ~w4485;
assign w4487 = ~w4479 & w4486;
assign w4488 = w4479 & ~w4486;
assign w4489 = ~w4487 & ~w4488;
assign w4490 = A_904 & A_905;
assign w4491 = (~w4490 & w4484) | (~w4490 & w13345) | (w4484 & w13345);
assign w4492 = A_901 & A_902;
assign w4493 = (~w4492 & w4477) | (~w4492 & w13346) | (w4477 & w13346);
assign w4494 = ~w4491 & w4493;
assign w4495 = w4491 & ~w4493;
assign w4496 = ~w4494 & ~w4495;
assign w4497 = ~w4479 & ~w4486;
assign w4498 = ~w4496 & w4497;
assign w4499 = ~w4491 & ~w4493;
assign w4500 = ~w4498 & ~w4499;
assign w4501 = w4497 & w4496;
assign w4502 = ~w4496 & ~w4497;
assign w4503 = ~w4501 & ~w4502;
assign w4504 = ~w4500 & ~w4503;
assign w4505 = ~w4489 & ~w4504;
assign w4506 = ~A_895 & A_896;
assign w4507 = A_895 & ~A_896;
assign w4508 = A_897 & ~w4507;
assign w4509 = ~w4506 & w4508;
assign w4510 = ~w4506 & ~w4507;
assign w4511 = ~A_897 & ~w4510;
assign w4512 = ~w4509 & ~w4511;
assign w4513 = ~A_898 & A_899;
assign w4514 = A_898 & ~A_899;
assign w4515 = A_900 & ~w4514;
assign w4516 = ~w4513 & w4515;
assign w4517 = ~w4513 & ~w4514;
assign w4518 = ~A_900 & ~w4517;
assign w4519 = ~w4516 & ~w4518;
assign w4520 = ~w4512 & w4519;
assign w4521 = w4512 & ~w4519;
assign w4522 = ~w4520 & ~w4521;
assign w4523 = A_898 & A_899;
assign w4524 = (~w4523 & w4517) | (~w4523 & w13347) | (w4517 & w13347);
assign w4525 = A_895 & A_896;
assign w4526 = (~w4525 & w4510) | (~w4525 & w13348) | (w4510 & w13348);
assign w4527 = ~w4524 & w4526;
assign w4528 = w4524 & ~w4526;
assign w4529 = ~w4527 & ~w4528;
assign w4530 = ~w4512 & ~w4519;
assign w4531 = ~w4529 & w4530;
assign w4532 = ~w4524 & ~w4526;
assign w4533 = ~w4531 & ~w4532;
assign w4534 = w4530 & w4529;
assign w4535 = ~w4529 & ~w4530;
assign w4536 = ~w4534 & ~w4535;
assign w4537 = ~w4533 & ~w4536;
assign w4538 = ~w4522 & ~w4537;
assign w4539 = ~w4505 & w4538;
assign w4540 = w4505 & ~w4538;
assign w4541 = ~w4539 & ~w4540;
assign w4542 = ~w4472 & w4541;
assign w4543 = w4472 & ~w4541;
assign w4544 = ~w4542 & ~w4543;
assign w4545 = ~w4403 & w4544;
assign w4546 = w4403 & ~w4544;
assign w4547 = ~w4545 & ~w4546;
assign w4548 = ~A_889 & A_890;
assign w4549 = A_889 & ~A_890;
assign w4550 = A_891 & ~w4549;
assign w4551 = ~w4548 & w4550;
assign w4552 = ~w4548 & ~w4549;
assign w4553 = ~A_891 & ~w4552;
assign w4554 = ~w4551 & ~w4553;
assign w4555 = ~A_892 & A_893;
assign w4556 = A_892 & ~A_893;
assign w4557 = A_894 & ~w4556;
assign w4558 = ~w4555 & w4557;
assign w4559 = ~w4555 & ~w4556;
assign w4560 = ~A_894 & ~w4559;
assign w4561 = ~w4558 & ~w4560;
assign w4562 = ~w4554 & w4561;
assign w4563 = w4554 & ~w4561;
assign w4564 = ~w4562 & ~w4563;
assign w4565 = A_892 & A_893;
assign w4566 = (~w4565 & w4559) | (~w4565 & w13349) | (w4559 & w13349);
assign w4567 = A_889 & A_890;
assign w4568 = (~w4567 & w4552) | (~w4567 & w13350) | (w4552 & w13350);
assign w4569 = ~w4566 & w4568;
assign w4570 = w4566 & ~w4568;
assign w4571 = ~w4569 & ~w4570;
assign w4572 = ~w4554 & ~w4561;
assign w4573 = ~w4571 & w4572;
assign w4574 = ~w4566 & ~w4568;
assign w4575 = ~w4573 & ~w4574;
assign w4576 = w4572 & w4571;
assign w4577 = ~w4571 & ~w4572;
assign w4578 = ~w4576 & ~w4577;
assign w4579 = ~w4575 & ~w4578;
assign w4580 = ~w4564 & ~w4579;
assign w4581 = ~A_883 & A_884;
assign w4582 = A_883 & ~A_884;
assign w4583 = A_885 & ~w4582;
assign w4584 = ~w4581 & w4583;
assign w4585 = ~w4581 & ~w4582;
assign w4586 = ~A_885 & ~w4585;
assign w4587 = ~w4584 & ~w4586;
assign w4588 = ~A_886 & A_887;
assign w4589 = A_886 & ~A_887;
assign w4590 = A_888 & ~w4589;
assign w4591 = ~w4588 & w4590;
assign w4592 = ~w4588 & ~w4589;
assign w4593 = ~A_888 & ~w4592;
assign w4594 = ~w4591 & ~w4593;
assign w4595 = ~w4587 & w4594;
assign w4596 = w4587 & ~w4594;
assign w4597 = ~w4595 & ~w4596;
assign w4598 = A_886 & A_887;
assign w4599 = (~w4598 & w4592) | (~w4598 & w13351) | (w4592 & w13351);
assign w4600 = A_883 & A_884;
assign w4601 = (~w4600 & w4585) | (~w4600 & w13352) | (w4585 & w13352);
assign w4602 = ~w4599 & w4601;
assign w4603 = w4599 & ~w4601;
assign w4604 = ~w4602 & ~w4603;
assign w4605 = ~w4587 & ~w4594;
assign w4606 = ~w4604 & w4605;
assign w4607 = ~w4599 & ~w4601;
assign w4608 = ~w4606 & ~w4607;
assign w4609 = w4605 & w4604;
assign w4610 = ~w4604 & ~w4605;
assign w4611 = ~w4609 & ~w4610;
assign w4612 = ~w4608 & ~w4611;
assign w4613 = ~w4597 & ~w4612;
assign w4614 = ~w4580 & w4613;
assign w4615 = w4580 & ~w4613;
assign w4616 = ~w4614 & ~w4615;
assign w4617 = ~A_877 & A_878;
assign w4618 = A_877 & ~A_878;
assign w4619 = A_879 & ~w4618;
assign w4620 = ~w4617 & w4619;
assign w4621 = ~w4617 & ~w4618;
assign w4622 = ~A_879 & ~w4621;
assign w4623 = ~w4620 & ~w4622;
assign w4624 = ~A_880 & A_881;
assign w4625 = A_880 & ~A_881;
assign w4626 = A_882 & ~w4625;
assign w4627 = ~w4624 & w4626;
assign w4628 = ~w4624 & ~w4625;
assign w4629 = ~A_882 & ~w4628;
assign w4630 = ~w4627 & ~w4629;
assign w4631 = ~w4623 & w4630;
assign w4632 = w4623 & ~w4630;
assign w4633 = ~w4631 & ~w4632;
assign w4634 = A_880 & A_881;
assign w4635 = (~w4634 & w4628) | (~w4634 & w13353) | (w4628 & w13353);
assign w4636 = A_877 & A_878;
assign w4637 = (~w4636 & w4621) | (~w4636 & w13354) | (w4621 & w13354);
assign w4638 = ~w4635 & w4637;
assign w4639 = w4635 & ~w4637;
assign w4640 = ~w4638 & ~w4639;
assign w4641 = ~w4623 & ~w4630;
assign w4642 = ~w4640 & w4641;
assign w4643 = ~w4635 & ~w4637;
assign w4644 = ~w4642 & ~w4643;
assign w4645 = w4641 & w4640;
assign w4646 = ~w4640 & ~w4641;
assign w4647 = ~w4645 & ~w4646;
assign w4648 = ~w4644 & ~w4647;
assign w4649 = ~w4633 & ~w4648;
assign w4650 = ~A_871 & A_872;
assign w4651 = A_871 & ~A_872;
assign w4652 = A_873 & ~w4651;
assign w4653 = ~w4650 & w4652;
assign w4654 = ~w4650 & ~w4651;
assign w4655 = ~A_873 & ~w4654;
assign w4656 = ~w4653 & ~w4655;
assign w4657 = ~A_874 & A_875;
assign w4658 = A_874 & ~A_875;
assign w4659 = A_876 & ~w4658;
assign w4660 = ~w4657 & w4659;
assign w4661 = ~w4657 & ~w4658;
assign w4662 = ~A_876 & ~w4661;
assign w4663 = ~w4660 & ~w4662;
assign w4664 = ~w4656 & w4663;
assign w4665 = w4656 & ~w4663;
assign w4666 = ~w4664 & ~w4665;
assign w4667 = A_874 & A_875;
assign w4668 = (~w4667 & w4661) | (~w4667 & w13355) | (w4661 & w13355);
assign w4669 = A_871 & A_872;
assign w4670 = (~w4669 & w4654) | (~w4669 & w13356) | (w4654 & w13356);
assign w4671 = ~w4668 & w4670;
assign w4672 = w4668 & ~w4670;
assign w4673 = ~w4671 & ~w4672;
assign w4674 = ~w4656 & ~w4663;
assign w4675 = ~w4673 & w4674;
assign w4676 = ~w4668 & ~w4670;
assign w4677 = ~w4675 & ~w4676;
assign w4678 = w4674 & w4673;
assign w4679 = ~w4673 & ~w4674;
assign w4680 = ~w4678 & ~w4679;
assign w4681 = ~w4677 & ~w4680;
assign w4682 = ~w4666 & ~w4681;
assign w4683 = ~w4649 & w4682;
assign w4684 = w4649 & ~w4682;
assign w4685 = ~w4683 & ~w4684;
assign w4686 = ~w4616 & w4685;
assign w4687 = w4616 & ~w4685;
assign w4688 = ~w4686 & ~w4687;
assign w4689 = ~A_865 & A_866;
assign w4690 = A_865 & ~A_866;
assign w4691 = A_867 & ~w4690;
assign w4692 = ~w4689 & w4691;
assign w4693 = ~w4689 & ~w4690;
assign w4694 = ~A_867 & ~w4693;
assign w4695 = ~w4692 & ~w4694;
assign w4696 = ~A_868 & A_869;
assign w4697 = A_868 & ~A_869;
assign w4698 = A_870 & ~w4697;
assign w4699 = ~w4696 & w4698;
assign w4700 = ~w4696 & ~w4697;
assign w4701 = ~A_870 & ~w4700;
assign w4702 = ~w4699 & ~w4701;
assign w4703 = ~w4695 & w4702;
assign w4704 = w4695 & ~w4702;
assign w4705 = ~w4703 & ~w4704;
assign w4706 = A_868 & A_869;
assign w4707 = (~w4706 & w4700) | (~w4706 & w13357) | (w4700 & w13357);
assign w4708 = A_865 & A_866;
assign w4709 = (~w4708 & w4693) | (~w4708 & w13358) | (w4693 & w13358);
assign w4710 = ~w4707 & w4709;
assign w4711 = w4707 & ~w4709;
assign w4712 = ~w4710 & ~w4711;
assign w4713 = ~w4695 & ~w4702;
assign w4714 = ~w4712 & w4713;
assign w4715 = ~w4707 & ~w4709;
assign w4716 = ~w4714 & ~w4715;
assign w4717 = w4713 & w4712;
assign w4718 = ~w4712 & ~w4713;
assign w4719 = ~w4717 & ~w4718;
assign w4720 = ~w4716 & ~w4719;
assign w4721 = ~w4705 & ~w4720;
assign w4722 = ~A_859 & A_860;
assign w4723 = A_859 & ~A_860;
assign w4724 = A_861 & ~w4723;
assign w4725 = ~w4722 & w4724;
assign w4726 = ~w4722 & ~w4723;
assign w4727 = ~A_861 & ~w4726;
assign w4728 = ~w4725 & ~w4727;
assign w4729 = ~A_862 & A_863;
assign w4730 = A_862 & ~A_863;
assign w4731 = A_864 & ~w4730;
assign w4732 = ~w4729 & w4731;
assign w4733 = ~w4729 & ~w4730;
assign w4734 = ~A_864 & ~w4733;
assign w4735 = ~w4732 & ~w4734;
assign w4736 = ~w4728 & w4735;
assign w4737 = w4728 & ~w4735;
assign w4738 = ~w4736 & ~w4737;
assign w4739 = A_862 & A_863;
assign w4740 = (~w4739 & w4733) | (~w4739 & w13359) | (w4733 & w13359);
assign w4741 = A_859 & A_860;
assign w4742 = (~w4741 & w4726) | (~w4741 & w13360) | (w4726 & w13360);
assign w4743 = ~w4740 & w4742;
assign w4744 = w4740 & ~w4742;
assign w4745 = ~w4743 & ~w4744;
assign w4746 = ~w4728 & ~w4735;
assign w4747 = ~w4745 & w4746;
assign w4748 = ~w4740 & ~w4742;
assign w4749 = ~w4747 & ~w4748;
assign w4750 = w4746 & w4745;
assign w4751 = ~w4745 & ~w4746;
assign w4752 = ~w4750 & ~w4751;
assign w4753 = ~w4749 & ~w4752;
assign w4754 = ~w4738 & ~w4753;
assign w4755 = ~w4721 & w4754;
assign w4756 = w4721 & ~w4754;
assign w4757 = ~w4755 & ~w4756;
assign w4758 = ~A_853 & A_854;
assign w4759 = A_853 & ~A_854;
assign w4760 = A_855 & ~w4759;
assign w4761 = ~w4758 & w4760;
assign w4762 = ~w4758 & ~w4759;
assign w4763 = ~A_855 & ~w4762;
assign w4764 = ~w4761 & ~w4763;
assign w4765 = ~A_856 & A_857;
assign w4766 = A_856 & ~A_857;
assign w4767 = A_858 & ~w4766;
assign w4768 = ~w4765 & w4767;
assign w4769 = ~w4765 & ~w4766;
assign w4770 = ~A_858 & ~w4769;
assign w4771 = ~w4768 & ~w4770;
assign w4772 = ~w4764 & w4771;
assign w4773 = w4764 & ~w4771;
assign w4774 = ~w4772 & ~w4773;
assign w4775 = A_856 & A_857;
assign w4776 = (~w4775 & w4769) | (~w4775 & w13361) | (w4769 & w13361);
assign w4777 = A_853 & A_854;
assign w4778 = (~w4777 & w4762) | (~w4777 & w13362) | (w4762 & w13362);
assign w4779 = ~w4776 & w4778;
assign w4780 = w4776 & ~w4778;
assign w4781 = ~w4779 & ~w4780;
assign w4782 = ~w4764 & ~w4771;
assign w4783 = ~w4781 & w4782;
assign w4784 = ~w4776 & ~w4778;
assign w4785 = ~w4783 & ~w4784;
assign w4786 = w4782 & w4781;
assign w4787 = ~w4781 & ~w4782;
assign w4788 = ~w4786 & ~w4787;
assign w4789 = ~w4785 & ~w4788;
assign w4790 = ~w4774 & ~w4789;
assign w4791 = ~A_847 & A_848;
assign w4792 = A_847 & ~A_848;
assign w4793 = A_849 & ~w4792;
assign w4794 = ~w4791 & w4793;
assign w4795 = ~w4791 & ~w4792;
assign w4796 = ~A_849 & ~w4795;
assign w4797 = ~w4794 & ~w4796;
assign w4798 = ~A_850 & A_851;
assign w4799 = A_850 & ~A_851;
assign w4800 = A_852 & ~w4799;
assign w4801 = ~w4798 & w4800;
assign w4802 = ~w4798 & ~w4799;
assign w4803 = ~A_852 & ~w4802;
assign w4804 = ~w4801 & ~w4803;
assign w4805 = ~w4797 & w4804;
assign w4806 = w4797 & ~w4804;
assign w4807 = ~w4805 & ~w4806;
assign w4808 = A_850 & A_851;
assign w4809 = (~w4808 & w4802) | (~w4808 & w13363) | (w4802 & w13363);
assign w4810 = A_847 & A_848;
assign w4811 = (~w4810 & w4795) | (~w4810 & w13364) | (w4795 & w13364);
assign w4812 = ~w4809 & w4811;
assign w4813 = w4809 & ~w4811;
assign w4814 = ~w4812 & ~w4813;
assign w4815 = ~w4797 & ~w4804;
assign w4816 = ~w4814 & w4815;
assign w4817 = ~w4809 & ~w4811;
assign w4818 = ~w4816 & ~w4817;
assign w4819 = w4815 & w4814;
assign w4820 = ~w4814 & ~w4815;
assign w4821 = ~w4819 & ~w4820;
assign w4822 = ~w4818 & ~w4821;
assign w4823 = ~w4807 & ~w4822;
assign w4824 = ~w4790 & w4823;
assign w4825 = w4790 & ~w4823;
assign w4826 = ~w4824 & ~w4825;
assign w4827 = ~w4757 & w4826;
assign w4828 = w4757 & ~w4826;
assign w4829 = ~w4827 & ~w4828;
assign w4830 = ~w4688 & w4829;
assign w4831 = w4688 & ~w4829;
assign w4832 = ~w4830 & ~w4831;
assign w4833 = ~w4547 & w4832;
assign w4834 = w4547 & ~w4832;
assign w4835 = ~w4833 & ~w4834;
assign w4836 = ~w4262 & ~w4835;
assign w4837 = ~w4258 & w4836;
assign w4838 = ~w4254 & w4837;
assign w4839 = ~w4254 & ~w4258;
assign w4840 = ~w4836 & ~w4839;
assign w4841 = ~w4838 & ~w4840;
assign w4842 = ~w4453 & ~w4464;
assign w4843 = ~w4467 & ~w4842;
assign w4844 = ~w4420 & ~w4453;
assign w4845 = ~w4435 & w4844;
assign w4846 = ~w4468 & w4845;
assign w4847 = ~w4420 & ~w4431;
assign w4848 = ~w4434 & ~w4847;
assign w4849 = ~w4846 & ~w4848;
assign w4850 = ~w4434 & w4844;
assign w4851 = ~w4435 & w4850;
assign w4852 = ~w4468 & ~w4847;
assign w4853 = w4851 & w4852;
assign w4854 = (w4843 & w4849) | (w4843 & w13847) | (w4849 & w13847);
assign w4855 = ~w4846 & w4848;
assign w4856 = w4846 & ~w4848;
assign w4857 = ~w4855 & ~w4856;
assign w4858 = ~w4843 & ~w4857;
assign w4859 = ~w4472 & ~w4541;
assign w4860 = ~w4858 & w13848;
assign w4861 = (~w4859 & w4858) | (~w4859 & w13849) | (w4858 & w13849);
assign w4862 = ~w4860 & ~w4861;
assign w4863 = ~w4522 & ~w4533;
assign w4864 = ~w4536 & ~w4863;
assign w4865 = ~w4489 & ~w4522;
assign w4866 = ~w4504 & w4865;
assign w4867 = ~w4537 & w4866;
assign w4868 = ~w4489 & ~w4500;
assign w4869 = ~w4503 & ~w4868;
assign w4870 = ~w4867 & w4869;
assign w4871 = w4867 & ~w4869;
assign w4872 = ~w4870 & ~w4871;
assign w4873 = ~w4864 & ~w4872;
assign w4874 = ~w4867 & ~w4869;
assign w4875 = ~w4503 & w4865;
assign w4876 = ~w4504 & w4875;
assign w4877 = ~w4537 & ~w4868;
assign w4878 = w4876 & w4877;
assign w4879 = (w4864 & w4874) | (w4864 & w13850) | (w4874 & w13850);
assign w4880 = ~w4873 & ~w4879;
assign w4881 = ~w4862 & w4880;
assign w4882 = ~w4858 & w13851;
assign w4883 = (w4859 & w4858) | (w4859 & w14059) | (w4858 & w14059);
assign w4884 = (~w4880 & w4883) | (~w4880 & w13852) | (w4883 & w13852);
assign w4885 = ~w4881 & ~w4884;
assign w4886 = ~w4381 & ~w4392;
assign w4887 = ~w4395 & ~w4886;
assign w4888 = ~w4348 & ~w4381;
assign w4889 = ~w4363 & w4888;
assign w4890 = ~w4396 & w4889;
assign w4891 = ~w4348 & ~w4359;
assign w4892 = ~w4362 & ~w4891;
assign w4893 = ~w4890 & w4892;
assign w4894 = w4890 & ~w4892;
assign w4895 = ~w4893 & ~w4894;
assign w4896 = ~w4887 & ~w4895;
assign w4897 = ~w4890 & ~w4892;
assign w4898 = ~w4362 & w4888;
assign w4899 = ~w4363 & w4898;
assign w4900 = ~w4396 & ~w4891;
assign w4901 = w4899 & w4900;
assign w4902 = (w4887 & w4897) | (w4887 & w13853) | (w4897 & w13853);
assign w4903 = ~w4896 & ~w4902;
assign w4904 = ~w4312 & ~w4323;
assign w4905 = ~w4326 & ~w4904;
assign w4906 = ~w4279 & ~w4312;
assign w4907 = ~w4294 & w4906;
assign w4908 = ~w4327 & w4907;
assign w4909 = ~w4279 & ~w4290;
assign w4910 = ~w4293 & ~w4909;
assign w4911 = ~w4908 & ~w4910;
assign w4912 = ~w4293 & w4906;
assign w4913 = ~w4294 & w4912;
assign w4914 = ~w4327 & ~w4909;
assign w4915 = w4913 & w4914;
assign w4916 = (w4905 & w4911) | (w4905 & w13529) | (w4911 & w13529);
assign w4917 = ~w4908 & w4910;
assign w4918 = w4908 & ~w4910;
assign w4919 = ~w4917 & ~w4918;
assign w4920 = ~w4905 & ~w4919;
assign w4921 = ~w4331 & ~w4400;
assign w4922 = ~w4920 & w13530;
assign w4923 = (w4921 & w4920) | (w4921 & w13531) | (w4920 & w13531);
assign w4924 = ~w4922 & ~w4923;
assign w4925 = ~w4903 & ~w4924;
assign w4926 = ~w4920 & w13532;
assign w4927 = (~w4921 & w4920) | (~w4921 & w13854) | (w4920 & w13854);
assign w4928 = (w4903 & w4927) | (w4903 & w13533) | (w4927 & w13533);
assign w4929 = ~w4403 & ~w4544;
assign w4930 = ~w4929 & ~w4928;
assign w4931 = ~w4925 & w4930;
assign w4932 = ~w4925 & ~w4928;
assign w4933 = w4929 & ~w4932;
assign w4934 = (~w4885 & w4933) | (~w4885 & w13855) | (w4933 & w13855);
assign w4935 = w4929 & ~w4928;
assign w4936 = ~w4925 & w4935;
assign w4937 = ~w4929 & ~w4932;
assign w4938 = ~w4936 & ~w4937;
assign w4939 = (w4885 & w4937) | (w4885 & w14060) | (w4937 & w14060);
assign w4940 = ~w4547 & ~w4832;
assign w4941 = (w4940 & w4938) | (w4940 & w13856) | (w4938 & w13856);
assign w4942 = ~w4934 & w4941;
assign w4943 = (~w4940 & w4939) | (~w4940 & w13857) | (w4939 & w13857);
assign w4944 = ~w4942 & ~w4943;
assign w4945 = ~w4666 & ~w4677;
assign w4946 = ~w4680 & ~w4945;
assign w4947 = ~w4633 & ~w4666;
assign w4948 = ~w4648 & w4947;
assign w4949 = ~w4681 & w4948;
assign w4950 = ~w4633 & ~w4644;
assign w4951 = ~w4647 & ~w4950;
assign w4952 = ~w4949 & w4951;
assign w4953 = w4949 & ~w4951;
assign w4954 = ~w4952 & ~w4953;
assign w4955 = ~w4946 & ~w4954;
assign w4956 = ~w4949 & ~w4951;
assign w4957 = ~w4647 & w4947;
assign w4958 = ~w4648 & w4957;
assign w4959 = ~w4681 & ~w4950;
assign w4960 = w4958 & w4959;
assign w4961 = (w4946 & w4956) | (w4946 & w13858) | (w4956 & w13858);
assign w4962 = ~w4955 & ~w4961;
assign w4963 = ~w4597 & ~w4608;
assign w4964 = ~w4611 & ~w4963;
assign w4965 = ~w4564 & ~w4597;
assign w4966 = ~w4579 & w4965;
assign w4967 = ~w4612 & w4966;
assign w4968 = ~w4564 & ~w4575;
assign w4969 = ~w4578 & ~w4968;
assign w4970 = ~w4967 & ~w4969;
assign w4971 = ~w4578 & w4965;
assign w4972 = ~w4579 & w4971;
assign w4973 = ~w4612 & ~w4968;
assign w4974 = w4972 & w4973;
assign w4975 = (w4964 & w4970) | (w4964 & w13534) | (w4970 & w13534);
assign w4976 = ~w4967 & w4969;
assign w4977 = w4967 & ~w4969;
assign w4978 = ~w4976 & ~w4977;
assign w4979 = ~w4964 & ~w4978;
assign w4980 = ~w4616 & ~w4685;
assign w4981 = ~w4979 & w13535;
assign w4982 = (w4980 & w4979) | (w4980 & w13859) | (w4979 & w13859);
assign w4983 = ~w4981 & ~w4982;
assign w4984 = ~w4962 & ~w4983;
assign w4985 = ~w4979 & w13536;
assign w4986 = (~w4980 & w4979) | (~w4980 & w13860) | (w4979 & w13860);
assign w4987 = (w4962 & w4986) | (w4962 & w13537) | (w4986 & w13537);
assign w4988 = ~w4688 & ~w4829;
assign w4989 = w4988 & ~w4987;
assign w4990 = ~w4984 & w4989;
assign w4991 = ~w4984 & ~w4987;
assign w4992 = ~w4988 & ~w4991;
assign w4993 = ~w4738 & ~w4749;
assign w4994 = ~w4752 & ~w4993;
assign w4995 = ~w4705 & ~w4738;
assign w4996 = ~w4720 & w4995;
assign w4997 = ~w4753 & w4996;
assign w4998 = ~w4705 & ~w4716;
assign w4999 = ~w4719 & ~w4998;
assign w5000 = ~w4997 & ~w4999;
assign w5001 = ~w4719 & w4995;
assign w5002 = ~w4720 & w5001;
assign w5003 = ~w4753 & ~w4998;
assign w5004 = w5002 & w5003;
assign w5005 = (w4994 & w5000) | (w4994 & w13861) | (w5000 & w13861);
assign w5006 = ~w4997 & w4999;
assign w5007 = w4997 & ~w4999;
assign w5008 = ~w5006 & ~w5007;
assign w5009 = ~w4994 & ~w5008;
assign w5010 = ~w4757 & ~w4826;
assign w5011 = ~w5009 & w13862;
assign w5012 = (~w5010 & w5009) | (~w5010 & w13863) | (w5009 & w13863);
assign w5013 = ~w5011 & ~w5012;
assign w5014 = ~w4807 & ~w4818;
assign w5015 = ~w4821 & ~w5014;
assign w5016 = ~w4774 & ~w4807;
assign w5017 = ~w4789 & w5016;
assign w5018 = ~w4822 & w5017;
assign w5019 = ~w4774 & ~w4785;
assign w5020 = ~w4788 & ~w5019;
assign w5021 = ~w5018 & w5020;
assign w5022 = w5018 & ~w5020;
assign w5023 = ~w5021 & ~w5022;
assign w5024 = ~w5015 & ~w5023;
assign w5025 = ~w5018 & ~w5020;
assign w5026 = ~w4788 & w5016;
assign w5027 = ~w4789 & w5026;
assign w5028 = ~w4822 & ~w5019;
assign w5029 = w5027 & w5028;
assign w5030 = (w5015 & w5025) | (w5015 & w13864) | (w5025 & w13864);
assign w5031 = ~w5024 & ~w5030;
assign w5032 = ~w5013 & w5031;
assign w5033 = ~w5009 & w13865;
assign w5034 = (w5010 & w5009) | (w5010 & w14061) | (w5009 & w14061);
assign w5035 = (~w5031 & w5034) | (~w5031 & w13866) | (w5034 & w13866);
assign w5036 = ~w5032 & ~w5035;
assign w5037 = (w5036 & w4992) | (w5036 & w13867) | (w4992 & w13867);
assign w5038 = ~w4988 & ~w4987;
assign w5039 = ~w4984 & w5038;
assign w5040 = w4988 & ~w4991;
assign w5041 = (~w5036 & w5040) | (~w5036 & w14062) | (w5040 & w14062);
assign w5042 = ~w5037 & ~w5041;
assign w5043 = ~w4944 & w5042;
assign w5044 = (~w4940 & w4938) | (~w4940 & w13868) | (w4938 & w13868);
assign w5045 = ~w4934 & w5044;
assign w5046 = (w4940 & w4939) | (w4940 & w13869) | (w4939 & w13869);
assign w5047 = ~w5045 & ~w5046;
assign w5048 = ~w5042 & ~w5047;
assign w5049 = ~w5043 & ~w5048;
assign w5050 = ~w4841 & w5049;
assign w5051 = ~w4258 & ~w4836;
assign w5052 = ~w4254 & w5051;
assign w5053 = w4836 & ~w4839;
assign w5054 = ~w5052 & ~w5053;
assign w5055 = ~w5049 & ~w5054;
assign w5056 = ~w5050 & ~w5055;
assign w5057 = A_202 & A_203;
assign w5058 = A_202 & ~A_203;
assign w5059 = ~A_202 & A_203;
assign w5060 = ~w5058 & ~w5059;
assign w5061 = (~w5057 & w5060) | (~w5057 & w12724) | (w5060 & w12724);
assign w5062 = A_199 & A_200;
assign w5063 = A_199 & ~A_200;
assign w5064 = ~A_199 & A_200;
assign w5065 = ~w5063 & ~w5064;
assign w5066 = (~w5062 & w5065) | (~w5062 & w12725) | (w5065 & w12725);
assign w5067 = w5061 & ~w5066;
assign w5068 = ~w5061 & w5066;
assign w5069 = A_201 & ~w5063;
assign w5070 = ~w5064 & w5069;
assign w5071 = ~A_201 & ~w5065;
assign w5072 = ~w5070 & ~w5071;
assign w5073 = A_204 & ~w5058;
assign w5074 = ~w5059 & w5073;
assign w5075 = ~A_204 & ~w5060;
assign w5076 = ~w5074 & ~w5075;
assign w5077 = ~w5072 & ~w5076;
assign w5078 = w5077 & w5079;
assign w5079 = ~w5067 & ~w5068;
assign w5080 = ~w5077 & ~w5079;
assign w5081 = ~w5078 & ~w5080;
assign w5082 = ~w5072 & w5076;
assign w5083 = w5072 & ~w5076;
assign w5084 = ~w5082 & ~w5083;
assign w5085 = w5077 & ~w5079;
assign w5086 = ~w5061 & ~w5066;
assign w5087 = ~w5085 & ~w5086;
assign w5088 = ~w5084 & ~w5087;
assign w5089 = ~w5081 & ~w5088;
assign w5090 = ~w5081 & ~w5087;
assign w5091 = A_208 & A_209;
assign w5092 = A_208 & ~A_209;
assign w5093 = ~A_208 & A_209;
assign w5094 = ~w5092 & ~w5093;
assign w5095 = (~w5091 & w5094) | (~w5091 & w12726) | (w5094 & w12726);
assign w5096 = A_205 & A_206;
assign w5097 = A_205 & ~A_206;
assign w5098 = ~A_205 & A_206;
assign w5099 = ~w5097 & ~w5098;
assign w5100 = (~w5096 & w5099) | (~w5096 & w12727) | (w5099 & w12727);
assign w5101 = ~w5095 & w5100;
assign w5102 = w5095 & ~w5100;
assign w5103 = ~w5101 & ~w5102;
assign w5104 = A_207 & ~w5097;
assign w5105 = ~w5098 & w5104;
assign w5106 = ~A_207 & ~w5099;
assign w5107 = ~w5105 & ~w5106;
assign w5108 = A_210 & ~w5092;
assign w5109 = ~w5093 & w5108;
assign w5110 = ~A_210 & ~w5094;
assign w5111 = ~w5109 & ~w5110;
assign w5112 = ~w5107 & ~w5111;
assign w5113 = ~w5103 & w5112;
assign w5114 = ~w5095 & ~w5100;
assign w5115 = ~w5113 & ~w5114;
assign w5116 = w5112 & w5103;
assign w5117 = ~w5103 & ~w5112;
assign w5118 = ~w5116 & ~w5117;
assign w5119 = ~w5115 & ~w5118;
assign w5120 = ~w5107 & w5111;
assign w5121 = w5107 & ~w5111;
assign w5122 = ~w5120 & ~w5121;
assign w5123 = ~w5084 & ~w5122;
assign w5124 = ~w5119 & w5123;
assign w5125 = ~w5090 & w5124;
assign w5126 = ~w5115 & ~w5122;
assign w5127 = ~w5118 & ~w5126;
assign w5128 = ~w5125 & w5127;
assign w5129 = w5125 & ~w5127;
assign w5130 = ~w5128 & ~w5129;
assign w5131 = ~w5089 & ~w5130;
assign w5132 = ~w5125 & ~w5127;
assign w5133 = ~w5118 & w5123;
assign w5134 = ~w5119 & w5133;
assign w5135 = ~w5090 & ~w5126;
assign w5136 = w5134 & w5135;
assign w5137 = (w5089 & w5132) | (w5089 & w13365) | (w5132 & w13365);
assign w5138 = ~w5131 & ~w5137;
assign w5139 = A_214 & A_215;
assign w5140 = A_214 & ~A_215;
assign w5141 = ~A_214 & A_215;
assign w5142 = ~w5140 & ~w5141;
assign w5143 = (~w5139 & w5142) | (~w5139 & w12728) | (w5142 & w12728);
assign w5144 = A_211 & A_212;
assign w5145 = A_211 & ~A_212;
assign w5146 = ~A_211 & A_212;
assign w5147 = ~w5145 & ~w5146;
assign w5148 = (~w5144 & w5147) | (~w5144 & w12729) | (w5147 & w12729);
assign w5149 = w5143 & ~w5148;
assign w5150 = ~w5143 & w5148;
assign w5151 = A_213 & ~w5145;
assign w5152 = ~w5146 & w5151;
assign w5153 = ~A_213 & ~w5147;
assign w5154 = ~w5152 & ~w5153;
assign w5155 = A_216 & ~w5140;
assign w5156 = ~w5141 & w5155;
assign w5157 = ~A_216 & ~w5142;
assign w5158 = ~w5156 & ~w5157;
assign w5159 = ~w5154 & ~w5158;
assign w5160 = w5159 & w5161;
assign w5161 = ~w5149 & ~w5150;
assign w5162 = ~w5159 & ~w5161;
assign w5163 = ~w5160 & ~w5162;
assign w5164 = ~w5154 & w5158;
assign w5165 = w5154 & ~w5158;
assign w5166 = ~w5164 & ~w5165;
assign w5167 = w5159 & ~w5161;
assign w5168 = ~w5143 & ~w5148;
assign w5169 = ~w5167 & ~w5168;
assign w5170 = ~w5166 & ~w5169;
assign w5171 = ~w5163 & ~w5170;
assign w5172 = ~w5163 & ~w5169;
assign w5173 = A_220 & A_221;
assign w5174 = A_220 & ~A_221;
assign w5175 = ~A_220 & A_221;
assign w5176 = ~w5174 & ~w5175;
assign w5177 = (~w5173 & w5176) | (~w5173 & w12730) | (w5176 & w12730);
assign w5178 = A_217 & A_218;
assign w5179 = A_217 & ~A_218;
assign w5180 = ~A_217 & A_218;
assign w5181 = ~w5179 & ~w5180;
assign w5182 = (~w5178 & w5181) | (~w5178 & w12731) | (w5181 & w12731);
assign w5183 = ~w5177 & w5182;
assign w5184 = w5177 & ~w5182;
assign w5185 = ~w5183 & ~w5184;
assign w5186 = A_219 & ~w5179;
assign w5187 = ~w5180 & w5186;
assign w5188 = ~A_219 & ~w5181;
assign w5189 = ~w5187 & ~w5188;
assign w5190 = A_222 & ~w5174;
assign w5191 = ~w5175 & w5190;
assign w5192 = ~A_222 & ~w5176;
assign w5193 = ~w5191 & ~w5192;
assign w5194 = ~w5189 & ~w5193;
assign w5195 = ~w5185 & w5194;
assign w5196 = ~w5177 & ~w5182;
assign w5197 = ~w5195 & ~w5196;
assign w5198 = w5194 & w5185;
assign w5199 = ~w5185 & ~w5194;
assign w5200 = ~w5198 & ~w5199;
assign w5201 = ~w5197 & ~w5200;
assign w5202 = ~w5189 & w5193;
assign w5203 = w5189 & ~w5193;
assign w5204 = ~w5202 & ~w5203;
assign w5205 = ~w5166 & ~w5204;
assign w5206 = ~w5201 & w5205;
assign w5207 = ~w5172 & w5206;
assign w5208 = ~w5197 & ~w5204;
assign w5209 = ~w5200 & ~w5208;
assign w5210 = ~w5207 & ~w5209;
assign w5211 = ~w5200 & w5205;
assign w5212 = ~w5201 & w5211;
assign w5213 = ~w5172 & ~w5208;
assign w5214 = w5212 & w5213;
assign w5215 = (w5171 & w5210) | (w5171 & w12984) | (w5210 & w12984);
assign w5216 = ~w5207 & w5209;
assign w5217 = w5207 & ~w5209;
assign w5218 = ~w5216 & ~w5217;
assign w5219 = ~w5171 & ~w5218;
assign w5220 = ~w5201 & ~w5204;
assign w5221 = ~w5166 & ~w5172;
assign w5222 = ~w5220 & w5221;
assign w5223 = w5220 & ~w5221;
assign w5224 = ~w5222 & ~w5223;
assign w5225 = ~w5119 & ~w5122;
assign w5226 = ~w5084 & ~w5090;
assign w5227 = ~w5225 & w5226;
assign w5228 = w5225 & ~w5226;
assign w5229 = ~w5227 & ~w5228;
assign w5230 = ~w5224 & ~w5229;
assign w5231 = ~w5219 & w12985;
assign w5232 = (w5230 & w5219) | (w5230 & w12986) | (w5219 & w12986);
assign w5233 = ~w5231 & ~w5232;
assign w5234 = ~w5138 & ~w5233;
assign w5235 = ~w5219 & w12987;
assign w5236 = (~w5230 & w5219) | (~w5230 & w13366) | (w5219 & w13366);
assign w5237 = (w5138 & w5236) | (w5138 & w12988) | (w5236 & w12988);
assign w5238 = ~w5224 & w5229;
assign w5239 = w5224 & ~w5229;
assign w5240 = ~w5238 & ~w5239;
assign w5241 = ~A_193 & A_194;
assign w5242 = A_193 & ~A_194;
assign w5243 = A_195 & ~w5242;
assign w5244 = ~w5241 & w5243;
assign w5245 = ~w5241 & ~w5242;
assign w5246 = ~A_195 & ~w5245;
assign w5247 = ~w5244 & ~w5246;
assign w5248 = ~A_196 & A_197;
assign w5249 = A_196 & ~A_197;
assign w5250 = A_198 & ~w5249;
assign w5251 = ~w5248 & w5250;
assign w5252 = ~w5248 & ~w5249;
assign w5253 = ~A_198 & ~w5252;
assign w5254 = ~w5251 & ~w5253;
assign w5255 = ~w5247 & w5254;
assign w5256 = w5247 & ~w5254;
assign w5257 = ~w5255 & ~w5256;
assign w5258 = A_196 & A_197;
assign w5259 = (~w5258 & w5252) | (~w5258 & w12732) | (w5252 & w12732);
assign w5260 = A_193 & A_194;
assign w5261 = (~w5260 & w5245) | (~w5260 & w12733) | (w5245 & w12733);
assign w5262 = ~w5259 & w5261;
assign w5263 = w5259 & ~w5261;
assign w5264 = ~w5262 & ~w5263;
assign w5265 = ~w5247 & ~w5254;
assign w5266 = ~w5264 & w5265;
assign w5267 = ~w5259 & ~w5261;
assign w5268 = ~w5266 & ~w5267;
assign w5269 = w5265 & w5264;
assign w5270 = ~w5264 & ~w5265;
assign w5271 = ~w5269 & ~w5270;
assign w5272 = ~w5268 & ~w5271;
assign w5273 = ~w5257 & ~w5272;
assign w5274 = ~A_187 & A_188;
assign w5275 = A_187 & ~A_188;
assign w5276 = A_189 & ~w5275;
assign w5277 = ~w5274 & w5276;
assign w5278 = ~w5274 & ~w5275;
assign w5279 = ~A_189 & ~w5278;
assign w5280 = ~w5277 & ~w5279;
assign w5281 = ~A_190 & A_191;
assign w5282 = A_190 & ~A_191;
assign w5283 = A_192 & ~w5282;
assign w5284 = ~w5281 & w5283;
assign w5285 = ~w5281 & ~w5282;
assign w5286 = ~A_192 & ~w5285;
assign w5287 = ~w5284 & ~w5286;
assign w5288 = ~w5280 & w5287;
assign w5289 = w5280 & ~w5287;
assign w5290 = ~w5288 & ~w5289;
assign w5291 = A_190 & A_191;
assign w5292 = (~w5291 & w5285) | (~w5291 & w12734) | (w5285 & w12734);
assign w5293 = A_187 & A_188;
assign w5294 = (~w5293 & w5278) | (~w5293 & w12735) | (w5278 & w12735);
assign w5295 = ~w5292 & w5294;
assign w5296 = w5292 & ~w5294;
assign w5297 = ~w5295 & ~w5296;
assign w5298 = ~w5280 & ~w5287;
assign w5299 = ~w5297 & w5298;
assign w5300 = ~w5292 & ~w5294;
assign w5301 = ~w5299 & ~w5300;
assign w5302 = w5298 & w5297;
assign w5303 = ~w5297 & ~w5298;
assign w5304 = ~w5302 & ~w5303;
assign w5305 = ~w5301 & ~w5304;
assign w5306 = ~w5290 & ~w5305;
assign w5307 = ~w5273 & w5306;
assign w5308 = w5273 & ~w5306;
assign w5309 = ~w5307 & ~w5308;
assign w5310 = ~A_181 & A_182;
assign w5311 = A_181 & ~A_182;
assign w5312 = A_183 & ~w5311;
assign w5313 = ~w5310 & w5312;
assign w5314 = ~w5310 & ~w5311;
assign w5315 = ~A_183 & ~w5314;
assign w5316 = ~w5313 & ~w5315;
assign w5317 = ~A_184 & A_185;
assign w5318 = A_184 & ~A_185;
assign w5319 = A_186 & ~w5318;
assign w5320 = ~w5317 & w5319;
assign w5321 = ~w5317 & ~w5318;
assign w5322 = ~A_186 & ~w5321;
assign w5323 = ~w5320 & ~w5322;
assign w5324 = ~w5316 & w5323;
assign w5325 = w5316 & ~w5323;
assign w5326 = ~w5324 & ~w5325;
assign w5327 = A_184 & A_185;
assign w5328 = (~w5327 & w5321) | (~w5327 & w12736) | (w5321 & w12736);
assign w5329 = A_181 & A_182;
assign w5330 = (~w5329 & w5314) | (~w5329 & w12737) | (w5314 & w12737);
assign w5331 = ~w5328 & w5330;
assign w5332 = w5328 & ~w5330;
assign w5333 = ~w5331 & ~w5332;
assign w5334 = ~w5316 & ~w5323;
assign w5335 = ~w5333 & w5334;
assign w5336 = ~w5328 & ~w5330;
assign w5337 = ~w5335 & ~w5336;
assign w5338 = w5334 & w5333;
assign w5339 = ~w5333 & ~w5334;
assign w5340 = ~w5338 & ~w5339;
assign w5341 = ~w5337 & ~w5340;
assign w5342 = ~w5326 & ~w5341;
assign w5343 = ~A_175 & A_176;
assign w5344 = A_175 & ~A_176;
assign w5345 = A_177 & ~w5344;
assign w5346 = ~w5343 & w5345;
assign w5347 = ~w5343 & ~w5344;
assign w5348 = ~A_177 & ~w5347;
assign w5349 = ~w5346 & ~w5348;
assign w5350 = ~A_178 & A_179;
assign w5351 = A_178 & ~A_179;
assign w5352 = A_180 & ~w5351;
assign w5353 = ~w5350 & w5352;
assign w5354 = ~w5350 & ~w5351;
assign w5355 = ~A_180 & ~w5354;
assign w5356 = ~w5353 & ~w5355;
assign w5357 = ~w5349 & w5356;
assign w5358 = w5349 & ~w5356;
assign w5359 = ~w5357 & ~w5358;
assign w5360 = A_178 & A_179;
assign w5361 = (~w5360 & w5354) | (~w5360 & w12738) | (w5354 & w12738);
assign w5362 = A_175 & A_176;
assign w5363 = (~w5362 & w5347) | (~w5362 & w12739) | (w5347 & w12739);
assign w5364 = ~w5361 & w5363;
assign w5365 = w5361 & ~w5363;
assign w5366 = ~w5364 & ~w5365;
assign w5367 = ~w5349 & ~w5356;
assign w5368 = ~w5366 & w5367;
assign w5369 = ~w5361 & ~w5363;
assign w5370 = ~w5368 & ~w5369;
assign w5371 = w5367 & w5366;
assign w5372 = ~w5366 & ~w5367;
assign w5373 = ~w5371 & ~w5372;
assign w5374 = ~w5370 & ~w5373;
assign w5375 = ~w5359 & ~w5374;
assign w5376 = ~w5342 & w5375;
assign w5377 = w5342 & ~w5375;
assign w5378 = ~w5376 & ~w5377;
assign w5379 = ~w5309 & w5378;
assign w5380 = w5309 & ~w5378;
assign w5381 = ~w5379 & ~w5380;
assign w5382 = ~w5240 & ~w5381;
assign w5383 = w5382 & ~w5237;
assign w5384 = ~w5234 & w5383;
assign w5385 = ~w5234 & ~w5237;
assign w5386 = ~w5382 & ~w5385;
assign w5387 = ~w5290 & ~w5301;
assign w5388 = ~w5304 & ~w5387;
assign w5389 = ~w5257 & ~w5290;
assign w5390 = ~w5272 & w5389;
assign w5391 = ~w5305 & w5390;
assign w5392 = ~w5257 & ~w5268;
assign w5393 = ~w5271 & ~w5392;
assign w5394 = ~w5391 & ~w5393;
assign w5395 = ~w5271 & w5389;
assign w5396 = ~w5272 & w5395;
assign w5397 = ~w5305 & ~w5392;
assign w5398 = w5396 & w5397;
assign w5399 = (w5388 & w5394) | (w5388 & w12989) | (w5394 & w12989);
assign w5400 = ~w5391 & w5393;
assign w5401 = w5391 & ~w5393;
assign w5402 = ~w5400 & ~w5401;
assign w5403 = ~w5388 & ~w5402;
assign w5404 = ~w5309 & ~w5378;
assign w5405 = ~w5403 & w13367;
assign w5406 = (~w5404 & w5403) | (~w5404 & w13368) | (w5403 & w13368);
assign w5407 = ~w5405 & ~w5406;
assign w5408 = ~w5359 & ~w5370;
assign w5409 = ~w5373 & ~w5408;
assign w5410 = ~w5326 & ~w5359;
assign w5411 = ~w5341 & w5410;
assign w5412 = ~w5374 & w5411;
assign w5413 = ~w5326 & ~w5337;
assign w5414 = ~w5340 & ~w5413;
assign w5415 = ~w5412 & w5414;
assign w5416 = w5412 & ~w5414;
assign w5417 = ~w5415 & ~w5416;
assign w5418 = ~w5409 & ~w5417;
assign w5419 = ~w5412 & ~w5414;
assign w5420 = ~w5340 & w5410;
assign w5421 = ~w5341 & w5420;
assign w5422 = ~w5374 & ~w5413;
assign w5423 = w5421 & w5422;
assign w5424 = (w5409 & w5419) | (w5409 & w13369) | (w5419 & w13369);
assign w5425 = ~w5418 & ~w5424;
assign w5426 = ~w5407 & w5425;
assign w5427 = ~w5403 & w12990;
assign w5428 = (w5404 & w5403) | (w5404 & w13370) | (w5403 & w13370);
assign w5429 = ~w5427 & ~w5428;
assign w5430 = ~w5425 & ~w5429;
assign w5431 = ~w5426 & ~w5430;
assign w5432 = (w5431 & w5386) | (w5431 & w13870) | (w5386 & w13870);
assign w5433 = ~w5382 & ~w5237;
assign w5434 = ~w5234 & w5433;
assign w5435 = w5382 & ~w5385;
assign w5436 = (~w5431 & w5435) | (~w5431 & w13871) | (w5435 & w13871);
assign w5437 = ~w5432 & ~w5436;
assign w5438 = A_238 & A_239;
assign w5439 = A_238 & ~A_239;
assign w5440 = ~A_238 & A_239;
assign w5441 = ~w5439 & ~w5440;
assign w5442 = (~w5438 & w5441) | (~w5438 & w12740) | (w5441 & w12740);
assign w5443 = A_235 & A_236;
assign w5444 = A_235 & ~A_236;
assign w5445 = ~A_235 & A_236;
assign w5446 = ~w5444 & ~w5445;
assign w5447 = (~w5443 & w5446) | (~w5443 & w12741) | (w5446 & w12741);
assign w5448 = w5442 & ~w5447;
assign w5449 = ~w5442 & w5447;
assign w5450 = A_237 & ~w5444;
assign w5451 = ~w5445 & w5450;
assign w5452 = ~A_237 & ~w5446;
assign w5453 = ~w5451 & ~w5452;
assign w5454 = A_240 & ~w5439;
assign w5455 = ~w5440 & w5454;
assign w5456 = ~A_240 & ~w5441;
assign w5457 = ~w5455 & ~w5456;
assign w5458 = ~w5453 & ~w5457;
assign w5459 = w5458 & w5460;
assign w5460 = ~w5448 & ~w5449;
assign w5461 = ~w5458 & ~w5460;
assign w5462 = ~w5459 & ~w5461;
assign w5463 = ~w5453 & w5457;
assign w5464 = w5453 & ~w5457;
assign w5465 = ~w5463 & ~w5464;
assign w5466 = w5458 & ~w5460;
assign w5467 = ~w5442 & ~w5447;
assign w5468 = ~w5466 & ~w5467;
assign w5469 = ~w5465 & ~w5468;
assign w5470 = ~w5462 & ~w5469;
assign w5471 = ~w5462 & ~w5468;
assign w5472 = A_244 & A_245;
assign w5473 = A_244 & ~A_245;
assign w5474 = ~A_244 & A_245;
assign w5475 = ~w5473 & ~w5474;
assign w5476 = (~w5472 & w5475) | (~w5472 & w12742) | (w5475 & w12742);
assign w5477 = A_241 & A_242;
assign w5478 = A_241 & ~A_242;
assign w5479 = ~A_241 & A_242;
assign w5480 = ~w5478 & ~w5479;
assign w5481 = (~w5477 & w5480) | (~w5477 & w12743) | (w5480 & w12743);
assign w5482 = ~w5476 & w5481;
assign w5483 = w5476 & ~w5481;
assign w5484 = ~w5482 & ~w5483;
assign w5485 = A_243 & ~w5478;
assign w5486 = ~w5479 & w5485;
assign w5487 = ~A_243 & ~w5480;
assign w5488 = ~w5486 & ~w5487;
assign w5489 = A_246 & ~w5473;
assign w5490 = ~w5474 & w5489;
assign w5491 = ~A_246 & ~w5475;
assign w5492 = ~w5490 & ~w5491;
assign w5493 = ~w5488 & ~w5492;
assign w5494 = ~w5484 & w5493;
assign w5495 = ~w5476 & ~w5481;
assign w5496 = ~w5494 & ~w5495;
assign w5497 = w5493 & w5484;
assign w5498 = ~w5484 & ~w5493;
assign w5499 = ~w5497 & ~w5498;
assign w5500 = ~w5496 & ~w5499;
assign w5501 = ~w5488 & w5492;
assign w5502 = w5488 & ~w5492;
assign w5503 = ~w5501 & ~w5502;
assign w5504 = ~w5465 & ~w5503;
assign w5505 = ~w5500 & w5504;
assign w5506 = ~w5471 & w5505;
assign w5507 = ~w5496 & ~w5503;
assign w5508 = ~w5499 & ~w5507;
assign w5509 = ~w5506 & ~w5508;
assign w5510 = ~w5499 & w5504;
assign w5511 = ~w5500 & w5510;
assign w5512 = ~w5471 & ~w5507;
assign w5513 = w5511 & w5512;
assign w5514 = (w5470 & w5509) | (w5470 & w12991) | (w5509 & w12991);
assign w5515 = ~w5506 & w5508;
assign w5516 = w5506 & ~w5508;
assign w5517 = ~w5515 & ~w5516;
assign w5518 = ~w5470 & ~w5517;
assign w5519 = ~w5500 & ~w5503;
assign w5520 = ~w5465 & ~w5471;
assign w5521 = ~w5519 & w5520;
assign w5522 = w5519 & ~w5520;
assign w5523 = ~w5521 & ~w5522;
assign w5524 = ~A_229 & A_230;
assign w5525 = A_229 & ~A_230;
assign w5526 = A_231 & ~w5525;
assign w5527 = ~w5524 & w5526;
assign w5528 = ~w5524 & ~w5525;
assign w5529 = ~A_231 & ~w5528;
assign w5530 = ~w5527 & ~w5529;
assign w5531 = ~A_232 & A_233;
assign w5532 = A_232 & ~A_233;
assign w5533 = A_234 & ~w5532;
assign w5534 = ~w5531 & w5533;
assign w5535 = ~w5531 & ~w5532;
assign w5536 = ~A_234 & ~w5535;
assign w5537 = ~w5534 & ~w5536;
assign w5538 = ~w5530 & w5537;
assign w5539 = w5530 & ~w5537;
assign w5540 = ~w5538 & ~w5539;
assign w5541 = A_232 & A_233;
assign w5542 = (~w5541 & w5535) | (~w5541 & w12744) | (w5535 & w12744);
assign w5543 = A_229 & A_230;
assign w5544 = (~w5543 & w5528) | (~w5543 & w12745) | (w5528 & w12745);
assign w5545 = ~w5542 & w5544;
assign w5546 = w5542 & ~w5544;
assign w5547 = ~w5545 & ~w5546;
assign w5548 = ~w5530 & ~w5537;
assign w5549 = ~w5547 & w5548;
assign w5550 = ~w5542 & ~w5544;
assign w5551 = ~w5549 & ~w5550;
assign w5552 = w5548 & w5547;
assign w5553 = ~w5547 & ~w5548;
assign w5554 = ~w5552 & ~w5553;
assign w5555 = ~w5551 & ~w5554;
assign w5556 = ~w5540 & ~w5555;
assign w5557 = ~A_223 & A_224;
assign w5558 = A_223 & ~A_224;
assign w5559 = A_225 & ~w5558;
assign w5560 = ~w5557 & w5559;
assign w5561 = ~w5557 & ~w5558;
assign w5562 = ~A_225 & ~w5561;
assign w5563 = ~w5560 & ~w5562;
assign w5564 = ~A_226 & A_227;
assign w5565 = A_226 & ~A_227;
assign w5566 = A_228 & ~w5565;
assign w5567 = ~w5564 & w5566;
assign w5568 = ~w5564 & ~w5565;
assign w5569 = ~A_228 & ~w5568;
assign w5570 = ~w5567 & ~w5569;
assign w5571 = ~w5563 & w5570;
assign w5572 = w5563 & ~w5570;
assign w5573 = ~w5571 & ~w5572;
assign w5574 = A_226 & A_227;
assign w5575 = (~w5574 & w5568) | (~w5574 & w12746) | (w5568 & w12746);
assign w5576 = A_223 & A_224;
assign w5577 = (~w5576 & w5561) | (~w5576 & w12747) | (w5561 & w12747);
assign w5578 = ~w5575 & w5577;
assign w5579 = w5575 & ~w5577;
assign w5580 = ~w5578 & ~w5579;
assign w5581 = ~w5563 & ~w5570;
assign w5582 = ~w5580 & w5581;
assign w5583 = ~w5575 & ~w5577;
assign w5584 = ~w5582 & ~w5583;
assign w5585 = w5581 & w5580;
assign w5586 = ~w5580 & ~w5581;
assign w5587 = ~w5585 & ~w5586;
assign w5588 = ~w5584 & ~w5587;
assign w5589 = ~w5573 & ~w5588;
assign w5590 = ~w5556 & w5589;
assign w5591 = w5556 & ~w5589;
assign w5592 = ~w5590 & ~w5591;
assign w5593 = ~w5523 & ~w5592;
assign w5594 = ~w5518 & w13371;
assign w5595 = (~w5593 & w5518) | (~w5593 & w13372) | (w5518 & w13372);
assign w5596 = ~w5594 & ~w5595;
assign w5597 = ~w5573 & ~w5584;
assign w5598 = ~w5587 & ~w5597;
assign w5599 = ~w5540 & ~w5573;
assign w5600 = ~w5555 & w5599;
assign w5601 = ~w5588 & w5600;
assign w5602 = ~w5540 & ~w5551;
assign w5603 = ~w5554 & ~w5602;
assign w5604 = ~w5601 & w5603;
assign w5605 = w5601 & ~w5603;
assign w5606 = ~w5604 & ~w5605;
assign w5607 = ~w5598 & ~w5606;
assign w5608 = ~w5601 & ~w5603;
assign w5609 = ~w5554 & w5599;
assign w5610 = ~w5555 & w5609;
assign w5611 = ~w5588 & ~w5602;
assign w5612 = w5610 & w5611;
assign w5613 = (w5598 & w5608) | (w5598 & w13373) | (w5608 & w13373);
assign w5614 = ~w5607 & ~w5613;
assign w5615 = ~w5596 & w5614;
assign w5616 = ~w5518 & w12992;
assign w5617 = (w5593 & w5518) | (w5593 & w13374) | (w5518 & w13374);
assign w5618 = ~w5616 & ~w5617;
assign w5619 = ~w5614 & ~w5618;
assign w5620 = ~w5615 & ~w5619;
assign w5621 = A_250 & A_251;
assign w5622 = A_250 & ~A_251;
assign w5623 = ~A_250 & A_251;
assign w5624 = ~w5622 & ~w5623;
assign w5625 = (~w5621 & w5624) | (~w5621 & w12748) | (w5624 & w12748);
assign w5626 = A_247 & A_248;
assign w5627 = A_247 & ~A_248;
assign w5628 = ~A_247 & A_248;
assign w5629 = ~w5627 & ~w5628;
assign w5630 = (~w5626 & w5629) | (~w5626 & w12749) | (w5629 & w12749);
assign w5631 = w5625 & ~w5630;
assign w5632 = ~w5625 & w5630;
assign w5633 = A_249 & ~w5627;
assign w5634 = ~w5628 & w5633;
assign w5635 = ~A_249 & ~w5629;
assign w5636 = ~w5634 & ~w5635;
assign w5637 = A_252 & ~w5622;
assign w5638 = ~w5623 & w5637;
assign w5639 = ~A_252 & ~w5624;
assign w5640 = ~w5638 & ~w5639;
assign w5641 = ~w5636 & ~w5640;
assign w5642 = w5641 & w5643;
assign w5643 = ~w5631 & ~w5632;
assign w5644 = ~w5641 & ~w5643;
assign w5645 = ~w5642 & ~w5644;
assign w5646 = ~w5636 & w5640;
assign w5647 = w5636 & ~w5640;
assign w5648 = ~w5646 & ~w5647;
assign w5649 = w5641 & ~w5643;
assign w5650 = ~w5625 & ~w5630;
assign w5651 = ~w5649 & ~w5650;
assign w5652 = ~w5648 & ~w5651;
assign w5653 = ~w5645 & ~w5652;
assign w5654 = ~w5645 & ~w5651;
assign w5655 = A_256 & A_257;
assign w5656 = A_256 & ~A_257;
assign w5657 = ~A_256 & A_257;
assign w5658 = ~w5656 & ~w5657;
assign w5659 = (~w5655 & w5658) | (~w5655 & w12750) | (w5658 & w12750);
assign w5660 = A_253 & A_254;
assign w5661 = A_253 & ~A_254;
assign w5662 = ~A_253 & A_254;
assign w5663 = ~w5661 & ~w5662;
assign w5664 = (~w5660 & w5663) | (~w5660 & w12751) | (w5663 & w12751);
assign w5665 = ~w5659 & w5664;
assign w5666 = w5659 & ~w5664;
assign w5667 = ~w5665 & ~w5666;
assign w5668 = A_255 & ~w5661;
assign w5669 = ~w5662 & w5668;
assign w5670 = ~A_255 & ~w5663;
assign w5671 = ~w5669 & ~w5670;
assign w5672 = A_258 & ~w5656;
assign w5673 = ~w5657 & w5672;
assign w5674 = ~A_258 & ~w5658;
assign w5675 = ~w5673 & ~w5674;
assign w5676 = ~w5671 & ~w5675;
assign w5677 = ~w5667 & w5676;
assign w5678 = ~w5659 & ~w5664;
assign w5679 = ~w5677 & ~w5678;
assign w5680 = w5676 & w5667;
assign w5681 = ~w5667 & ~w5676;
assign w5682 = ~w5680 & ~w5681;
assign w5683 = ~w5679 & ~w5682;
assign w5684 = ~w5671 & w5675;
assign w5685 = w5671 & ~w5675;
assign w5686 = ~w5684 & ~w5685;
assign w5687 = ~w5648 & ~w5686;
assign w5688 = ~w5683 & w5687;
assign w5689 = ~w5654 & w5688;
assign w5690 = ~w5679 & ~w5686;
assign w5691 = ~w5682 & ~w5690;
assign w5692 = ~w5689 & w5691;
assign w5693 = w5689 & ~w5691;
assign w5694 = ~w5692 & ~w5693;
assign w5695 = ~w5653 & ~w5694;
assign w5696 = ~w5689 & ~w5691;
assign w5697 = ~w5682 & w5687;
assign w5698 = ~w5683 & w5697;
assign w5699 = ~w5654 & ~w5690;
assign w5700 = w5698 & w5699;
assign w5701 = (w5653 & w5696) | (w5653 & w13375) | (w5696 & w13375);
assign w5702 = ~w5695 & ~w5701;
assign w5703 = A_262 & A_263;
assign w5704 = A_262 & ~A_263;
assign w5705 = ~A_262 & A_263;
assign w5706 = ~w5704 & ~w5705;
assign w5707 = (~w5703 & w5706) | (~w5703 & w12752) | (w5706 & w12752);
assign w5708 = A_259 & A_260;
assign w5709 = A_259 & ~A_260;
assign w5710 = ~A_259 & A_260;
assign w5711 = ~w5709 & ~w5710;
assign w5712 = (~w5708 & w5711) | (~w5708 & w12753) | (w5711 & w12753);
assign w5713 = w5707 & ~w5712;
assign w5714 = ~w5707 & w5712;
assign w5715 = A_261 & ~w5709;
assign w5716 = ~w5710 & w5715;
assign w5717 = ~A_261 & ~w5711;
assign w5718 = ~w5716 & ~w5717;
assign w5719 = A_264 & ~w5704;
assign w5720 = ~w5705 & w5719;
assign w5721 = ~A_264 & ~w5706;
assign w5722 = ~w5720 & ~w5721;
assign w5723 = ~w5718 & ~w5722;
assign w5724 = w5723 & w5725;
assign w5725 = ~w5713 & ~w5714;
assign w5726 = ~w5723 & ~w5725;
assign w5727 = ~w5724 & ~w5726;
assign w5728 = ~w5718 & w5722;
assign w5729 = w5718 & ~w5722;
assign w5730 = ~w5728 & ~w5729;
assign w5731 = w5723 & ~w5725;
assign w5732 = ~w5707 & ~w5712;
assign w5733 = ~w5731 & ~w5732;
assign w5734 = ~w5730 & ~w5733;
assign w5735 = ~w5727 & ~w5734;
assign w5736 = ~w5727 & ~w5733;
assign w5737 = A_268 & A_269;
assign w5738 = A_268 & ~A_269;
assign w5739 = ~A_268 & A_269;
assign w5740 = ~w5738 & ~w5739;
assign w5741 = (~w5737 & w5740) | (~w5737 & w12754) | (w5740 & w12754);
assign w5742 = A_265 & A_266;
assign w5743 = A_265 & ~A_266;
assign w5744 = ~A_265 & A_266;
assign w5745 = ~w5743 & ~w5744;
assign w5746 = (~w5742 & w5745) | (~w5742 & w12755) | (w5745 & w12755);
assign w5747 = ~w5741 & w5746;
assign w5748 = w5741 & ~w5746;
assign w5749 = ~w5747 & ~w5748;
assign w5750 = A_267 & ~w5743;
assign w5751 = ~w5744 & w5750;
assign w5752 = ~A_267 & ~w5745;
assign w5753 = ~w5751 & ~w5752;
assign w5754 = A_270 & ~w5738;
assign w5755 = ~w5739 & w5754;
assign w5756 = ~A_270 & ~w5740;
assign w5757 = ~w5755 & ~w5756;
assign w5758 = ~w5753 & ~w5757;
assign w5759 = ~w5749 & w5758;
assign w5760 = ~w5741 & ~w5746;
assign w5761 = ~w5759 & ~w5760;
assign w5762 = w5758 & w5749;
assign w5763 = ~w5749 & ~w5758;
assign w5764 = ~w5762 & ~w5763;
assign w5765 = ~w5761 & ~w5764;
assign w5766 = ~w5753 & w5757;
assign w5767 = w5753 & ~w5757;
assign w5768 = ~w5766 & ~w5767;
assign w5769 = ~w5730 & ~w5768;
assign w5770 = ~w5765 & w5769;
assign w5771 = ~w5736 & w5770;
assign w5772 = ~w5761 & ~w5768;
assign w5773 = ~w5764 & ~w5772;
assign w5774 = ~w5771 & ~w5773;
assign w5775 = ~w5764 & w5769;
assign w5776 = ~w5765 & w5775;
assign w5777 = ~w5736 & ~w5772;
assign w5778 = w5776 & w5777;
assign w5779 = (w5735 & w5774) | (w5735 & w12993) | (w5774 & w12993);
assign w5780 = ~w5771 & w5773;
assign w5781 = w5771 & ~w5773;
assign w5782 = ~w5780 & ~w5781;
assign w5783 = ~w5735 & ~w5782;
assign w5784 = ~w5765 & ~w5768;
assign w5785 = ~w5730 & ~w5736;
assign w5786 = ~w5784 & w5785;
assign w5787 = w5784 & ~w5785;
assign w5788 = ~w5786 & ~w5787;
assign w5789 = ~w5683 & ~w5686;
assign w5790 = ~w5648 & ~w5654;
assign w5791 = ~w5789 & w5790;
assign w5792 = w5789 & ~w5790;
assign w5793 = ~w5791 & ~w5792;
assign w5794 = ~w5788 & ~w5793;
assign w5795 = ~w5783 & w12994;
assign w5796 = (w5794 & w5783) | (w5794 & w12995) | (w5783 & w12995);
assign w5797 = ~w5795 & ~w5796;
assign w5798 = ~w5702 & ~w5797;
assign w5799 = ~w5783 & w12996;
assign w5800 = (~w5794 & w5783) | (~w5794 & w13376) | (w5783 & w13376);
assign w5801 = (w5702 & w5800) | (w5702 & w12997) | (w5800 & w12997);
assign w5802 = ~w5788 & w5793;
assign w5803 = w5788 & ~w5793;
assign w5804 = ~w5802 & ~w5803;
assign w5805 = ~w5523 & w5592;
assign w5806 = w5523 & ~w5592;
assign w5807 = ~w5805 & ~w5806;
assign w5808 = ~w5804 & ~w5807;
assign w5809 = ~w5808 & ~w5801;
assign w5810 = ~w5798 & w5809;
assign w5811 = ~w5798 & ~w5801;
assign w5812 = w5808 & ~w5811;
assign w5813 = (~w5620 & w5812) | (~w5620 & w13377) | (w5812 & w13377);
assign w5814 = w5808 & ~w5801;
assign w5815 = ~w5798 & w5814;
assign w5816 = ~w5808 & ~w5811;
assign w5817 = ~w5815 & ~w5816;
assign w5818 = (w5620 & w5816) | (w5620 & w13872) | (w5816 & w13872);
assign w5819 = ~w5804 & w5807;
assign w5820 = w5804 & ~w5807;
assign w5821 = ~w5819 & ~w5820;
assign w5822 = ~w5240 & w5381;
assign w5823 = w5240 & ~w5381;
assign w5824 = ~w5822 & ~w5823;
assign w5825 = ~w5821 & ~w5824;
assign w5826 = (~w5825 & w5817) | (~w5825 & w13378) | (w5817 & w13378);
assign w5827 = ~w5813 & w5826;
assign w5828 = (w5825 & w5818) | (w5825 & w13379) | (w5818 & w13379);
assign w5829 = ~w5827 & ~w5828;
assign w5830 = ~w5437 & ~w5829;
assign w5831 = (w5825 & w5817) | (w5825 & w13380) | (w5817 & w13380);
assign w5832 = ~w5813 & w5831;
assign w5833 = (~w5825 & w5818) | (~w5825 & w13381) | (w5818 & w13381);
assign w5834 = ~w5832 & ~w5833;
assign w5835 = w5437 & ~w5834;
assign w5836 = ~w5821 & w5824;
assign w5837 = w5821 & ~w5824;
assign w5838 = ~w5836 & ~w5837;
assign w5839 = ~A_169 & A_170;
assign w5840 = A_169 & ~A_170;
assign w5841 = A_171 & ~w5840;
assign w5842 = ~w5839 & w5841;
assign w5843 = ~w5839 & ~w5840;
assign w5844 = ~A_171 & ~w5843;
assign w5845 = ~w5842 & ~w5844;
assign w5846 = ~A_172 & A_173;
assign w5847 = A_172 & ~A_173;
assign w5848 = A_174 & ~w5847;
assign w5849 = ~w5846 & w5848;
assign w5850 = ~w5846 & ~w5847;
assign w5851 = ~A_174 & ~w5850;
assign w5852 = ~w5849 & ~w5851;
assign w5853 = ~w5845 & w5852;
assign w5854 = w5845 & ~w5852;
assign w5855 = ~w5853 & ~w5854;
assign w5856 = A_172 & A_173;
assign w5857 = (~w5856 & w5850) | (~w5856 & w12756) | (w5850 & w12756);
assign w5858 = A_169 & A_170;
assign w5859 = (~w5858 & w5843) | (~w5858 & w12757) | (w5843 & w12757);
assign w5860 = ~w5857 & w5859;
assign w5861 = w5857 & ~w5859;
assign w5862 = ~w5860 & ~w5861;
assign w5863 = ~w5845 & ~w5852;
assign w5864 = ~w5862 & w5863;
assign w5865 = ~w5857 & ~w5859;
assign w5866 = ~w5864 & ~w5865;
assign w5867 = w5863 & w5862;
assign w5868 = ~w5862 & ~w5863;
assign w5869 = ~w5867 & ~w5868;
assign w5870 = ~w5866 & ~w5869;
assign w5871 = ~w5855 & ~w5870;
assign w5872 = ~A_163 & A_164;
assign w5873 = A_163 & ~A_164;
assign w5874 = A_165 & ~w5873;
assign w5875 = ~w5872 & w5874;
assign w5876 = ~w5872 & ~w5873;
assign w5877 = ~A_165 & ~w5876;
assign w5878 = ~w5875 & ~w5877;
assign w5879 = ~A_166 & A_167;
assign w5880 = A_166 & ~A_167;
assign w5881 = A_168 & ~w5880;
assign w5882 = ~w5879 & w5881;
assign w5883 = ~w5879 & ~w5880;
assign w5884 = ~A_168 & ~w5883;
assign w5885 = ~w5882 & ~w5884;
assign w5886 = ~w5878 & w5885;
assign w5887 = w5878 & ~w5885;
assign w5888 = ~w5886 & ~w5887;
assign w5889 = A_166 & A_167;
assign w5890 = (~w5889 & w5883) | (~w5889 & w12758) | (w5883 & w12758);
assign w5891 = A_163 & A_164;
assign w5892 = (~w5891 & w5876) | (~w5891 & w12759) | (w5876 & w12759);
assign w5893 = ~w5890 & w5892;
assign w5894 = w5890 & ~w5892;
assign w5895 = ~w5893 & ~w5894;
assign w5896 = ~w5878 & ~w5885;
assign w5897 = ~w5895 & w5896;
assign w5898 = ~w5890 & ~w5892;
assign w5899 = ~w5897 & ~w5898;
assign w5900 = w5896 & w5895;
assign w5901 = ~w5895 & ~w5896;
assign w5902 = ~w5900 & ~w5901;
assign w5903 = ~w5899 & ~w5902;
assign w5904 = ~w5888 & ~w5903;
assign w5905 = ~w5871 & w5904;
assign w5906 = w5871 & ~w5904;
assign w5907 = ~w5905 & ~w5906;
assign w5908 = ~A_157 & A_158;
assign w5909 = A_157 & ~A_158;
assign w5910 = A_159 & ~w5909;
assign w5911 = ~w5908 & w5910;
assign w5912 = ~w5908 & ~w5909;
assign w5913 = ~A_159 & ~w5912;
assign w5914 = ~w5911 & ~w5913;
assign w5915 = ~A_160 & A_161;
assign w5916 = A_160 & ~A_161;
assign w5917 = A_162 & ~w5916;
assign w5918 = ~w5915 & w5917;
assign w5919 = ~w5915 & ~w5916;
assign w5920 = ~A_162 & ~w5919;
assign w5921 = ~w5918 & ~w5920;
assign w5922 = ~w5914 & w5921;
assign w5923 = w5914 & ~w5921;
assign w5924 = ~w5922 & ~w5923;
assign w5925 = A_160 & A_161;
assign w5926 = (~w5925 & w5919) | (~w5925 & w12760) | (w5919 & w12760);
assign w5927 = A_157 & A_158;
assign w5928 = (~w5927 & w5912) | (~w5927 & w12761) | (w5912 & w12761);
assign w5929 = ~w5926 & w5928;
assign w5930 = w5926 & ~w5928;
assign w5931 = ~w5929 & ~w5930;
assign w5932 = ~w5914 & ~w5921;
assign w5933 = ~w5931 & w5932;
assign w5934 = ~w5926 & ~w5928;
assign w5935 = ~w5933 & ~w5934;
assign w5936 = w5932 & w5931;
assign w5937 = ~w5931 & ~w5932;
assign w5938 = ~w5936 & ~w5937;
assign w5939 = ~w5935 & ~w5938;
assign w5940 = ~w5924 & ~w5939;
assign w5941 = ~A_151 & A_152;
assign w5942 = A_151 & ~A_152;
assign w5943 = A_153 & ~w5942;
assign w5944 = ~w5941 & w5943;
assign w5945 = ~w5941 & ~w5942;
assign w5946 = ~A_153 & ~w5945;
assign w5947 = ~w5944 & ~w5946;
assign w5948 = ~A_154 & A_155;
assign w5949 = A_154 & ~A_155;
assign w5950 = A_156 & ~w5949;
assign w5951 = ~w5948 & w5950;
assign w5952 = ~w5948 & ~w5949;
assign w5953 = ~A_156 & ~w5952;
assign w5954 = ~w5951 & ~w5953;
assign w5955 = ~w5947 & w5954;
assign w5956 = w5947 & ~w5954;
assign w5957 = ~w5955 & ~w5956;
assign w5958 = A_154 & A_155;
assign w5959 = (~w5958 & w5952) | (~w5958 & w12762) | (w5952 & w12762);
assign w5960 = A_151 & A_152;
assign w5961 = (~w5960 & w5945) | (~w5960 & w12763) | (w5945 & w12763);
assign w5962 = ~w5959 & w5961;
assign w5963 = w5959 & ~w5961;
assign w5964 = ~w5962 & ~w5963;
assign w5965 = ~w5947 & ~w5954;
assign w5966 = ~w5964 & w5965;
assign w5967 = ~w5959 & ~w5961;
assign w5968 = ~w5966 & ~w5967;
assign w5969 = w5965 & w5964;
assign w5970 = ~w5964 & ~w5965;
assign w5971 = ~w5969 & ~w5970;
assign w5972 = ~w5968 & ~w5971;
assign w5973 = ~w5957 & ~w5972;
assign w5974 = ~w5940 & w5973;
assign w5975 = w5940 & ~w5973;
assign w5976 = ~w5974 & ~w5975;
assign w5977 = ~w5907 & w5976;
assign w5978 = w5907 & ~w5976;
assign w5979 = ~w5977 & ~w5978;
assign w5980 = ~A_145 & A_146;
assign w5981 = A_145 & ~A_146;
assign w5982 = A_147 & ~w5981;
assign w5983 = ~w5980 & w5982;
assign w5984 = ~w5980 & ~w5981;
assign w5985 = ~A_147 & ~w5984;
assign w5986 = ~w5983 & ~w5985;
assign w5987 = ~A_148 & A_149;
assign w5988 = A_148 & ~A_149;
assign w5989 = A_150 & ~w5988;
assign w5990 = ~w5987 & w5989;
assign w5991 = ~w5987 & ~w5988;
assign w5992 = ~A_150 & ~w5991;
assign w5993 = ~w5990 & ~w5992;
assign w5994 = ~w5986 & w5993;
assign w5995 = w5986 & ~w5993;
assign w5996 = ~w5994 & ~w5995;
assign w5997 = A_148 & A_149;
assign w5998 = (~w5997 & w5991) | (~w5997 & w12764) | (w5991 & w12764);
assign w5999 = A_145 & A_146;
assign w6000 = (~w5999 & w5984) | (~w5999 & w12765) | (w5984 & w12765);
assign w6001 = ~w5998 & w6000;
assign w6002 = w5998 & ~w6000;
assign w6003 = ~w6001 & ~w6002;
assign w6004 = ~w5986 & ~w5993;
assign w6005 = ~w6003 & w6004;
assign w6006 = ~w5998 & ~w6000;
assign w6007 = ~w6005 & ~w6006;
assign w6008 = w6004 & w6003;
assign w6009 = ~w6003 & ~w6004;
assign w6010 = ~w6008 & ~w6009;
assign w6011 = ~w6007 & ~w6010;
assign w6012 = ~w5996 & ~w6011;
assign w6013 = ~A_139 & A_140;
assign w6014 = A_139 & ~A_140;
assign w6015 = A_141 & ~w6014;
assign w6016 = ~w6013 & w6015;
assign w6017 = ~w6013 & ~w6014;
assign w6018 = ~A_141 & ~w6017;
assign w6019 = ~w6016 & ~w6018;
assign w6020 = ~A_142 & A_143;
assign w6021 = A_142 & ~A_143;
assign w6022 = A_144 & ~w6021;
assign w6023 = ~w6020 & w6022;
assign w6024 = ~w6020 & ~w6021;
assign w6025 = ~A_144 & ~w6024;
assign w6026 = ~w6023 & ~w6025;
assign w6027 = ~w6019 & w6026;
assign w6028 = w6019 & ~w6026;
assign w6029 = ~w6027 & ~w6028;
assign w6030 = A_142 & A_143;
assign w6031 = (~w6030 & w6024) | (~w6030 & w12766) | (w6024 & w12766);
assign w6032 = A_139 & A_140;
assign w6033 = (~w6032 & w6017) | (~w6032 & w12767) | (w6017 & w12767);
assign w6034 = ~w6031 & w6033;
assign w6035 = w6031 & ~w6033;
assign w6036 = ~w6034 & ~w6035;
assign w6037 = ~w6019 & ~w6026;
assign w6038 = ~w6036 & w6037;
assign w6039 = ~w6031 & ~w6033;
assign w6040 = ~w6038 & ~w6039;
assign w6041 = w6037 & w6036;
assign w6042 = ~w6036 & ~w6037;
assign w6043 = ~w6041 & ~w6042;
assign w6044 = ~w6040 & ~w6043;
assign w6045 = ~w6029 & ~w6044;
assign w6046 = ~w6012 & w6045;
assign w6047 = w6012 & ~w6045;
assign w6048 = ~w6046 & ~w6047;
assign w6049 = ~A_133 & A_134;
assign w6050 = A_133 & ~A_134;
assign w6051 = A_135 & ~w6050;
assign w6052 = ~w6049 & w6051;
assign w6053 = ~w6049 & ~w6050;
assign w6054 = ~A_135 & ~w6053;
assign w6055 = ~w6052 & ~w6054;
assign w6056 = ~A_136 & A_137;
assign w6057 = A_136 & ~A_137;
assign w6058 = A_138 & ~w6057;
assign w6059 = ~w6056 & w6058;
assign w6060 = ~w6056 & ~w6057;
assign w6061 = ~A_138 & ~w6060;
assign w6062 = ~w6059 & ~w6061;
assign w6063 = ~w6055 & w6062;
assign w6064 = w6055 & ~w6062;
assign w6065 = ~w6063 & ~w6064;
assign w6066 = A_136 & A_137;
assign w6067 = (~w6066 & w6060) | (~w6066 & w12768) | (w6060 & w12768);
assign w6068 = A_133 & A_134;
assign w6069 = (~w6068 & w6053) | (~w6068 & w12769) | (w6053 & w12769);
assign w6070 = ~w6067 & w6069;
assign w6071 = w6067 & ~w6069;
assign w6072 = ~w6070 & ~w6071;
assign w6073 = ~w6055 & ~w6062;
assign w6074 = ~w6072 & w6073;
assign w6075 = ~w6067 & ~w6069;
assign w6076 = ~w6074 & ~w6075;
assign w6077 = w6073 & w6072;
assign w6078 = ~w6072 & ~w6073;
assign w6079 = ~w6077 & ~w6078;
assign w6080 = ~w6076 & ~w6079;
assign w6081 = ~w6065 & ~w6080;
assign w6082 = ~A_127 & A_128;
assign w6083 = A_127 & ~A_128;
assign w6084 = A_129 & ~w6083;
assign w6085 = ~w6082 & w6084;
assign w6086 = ~w6082 & ~w6083;
assign w6087 = ~A_129 & ~w6086;
assign w6088 = ~w6085 & ~w6087;
assign w6089 = ~A_130 & A_131;
assign w6090 = A_130 & ~A_131;
assign w6091 = A_132 & ~w6090;
assign w6092 = ~w6089 & w6091;
assign w6093 = ~w6089 & ~w6090;
assign w6094 = ~A_132 & ~w6093;
assign w6095 = ~w6092 & ~w6094;
assign w6096 = ~w6088 & w6095;
assign w6097 = w6088 & ~w6095;
assign w6098 = ~w6096 & ~w6097;
assign w6099 = A_130 & A_131;
assign w6100 = (~w6099 & w6093) | (~w6099 & w12770) | (w6093 & w12770);
assign w6101 = A_127 & A_128;
assign w6102 = (~w6101 & w6086) | (~w6101 & w12771) | (w6086 & w12771);
assign w6103 = ~w6100 & w6102;
assign w6104 = w6100 & ~w6102;
assign w6105 = ~w6103 & ~w6104;
assign w6106 = ~w6088 & ~w6095;
assign w6107 = ~w6105 & w6106;
assign w6108 = ~w6100 & ~w6102;
assign w6109 = ~w6107 & ~w6108;
assign w6110 = w6106 & w6105;
assign w6111 = ~w6105 & ~w6106;
assign w6112 = ~w6110 & ~w6111;
assign w6113 = ~w6109 & ~w6112;
assign w6114 = ~w6098 & ~w6113;
assign w6115 = ~w6081 & w6114;
assign w6116 = w6081 & ~w6114;
assign w6117 = ~w6115 & ~w6116;
assign w6118 = ~w6048 & w6117;
assign w6119 = w6048 & ~w6117;
assign w6120 = ~w6118 & ~w6119;
assign w6121 = ~w5979 & w6120;
assign w6122 = w5979 & ~w6120;
assign w6123 = ~w6121 & ~w6122;
assign w6124 = ~A_121 & A_122;
assign w6125 = A_121 & ~A_122;
assign w6126 = A_123 & ~w6125;
assign w6127 = ~w6124 & w6126;
assign w6128 = ~w6124 & ~w6125;
assign w6129 = ~A_123 & ~w6128;
assign w6130 = ~w6127 & ~w6129;
assign w6131 = ~A_124 & A_125;
assign w6132 = A_124 & ~A_125;
assign w6133 = A_126 & ~w6132;
assign w6134 = ~w6131 & w6133;
assign w6135 = ~w6131 & ~w6132;
assign w6136 = ~A_126 & ~w6135;
assign w6137 = ~w6134 & ~w6136;
assign w6138 = ~w6130 & w6137;
assign w6139 = w6130 & ~w6137;
assign w6140 = ~w6138 & ~w6139;
assign w6141 = A_124 & A_125;
assign w6142 = (~w6141 & w6135) | (~w6141 & w12772) | (w6135 & w12772);
assign w6143 = A_121 & A_122;
assign w6144 = (~w6143 & w6128) | (~w6143 & w12773) | (w6128 & w12773);
assign w6145 = ~w6142 & w6144;
assign w6146 = w6142 & ~w6144;
assign w6147 = ~w6145 & ~w6146;
assign w6148 = ~w6130 & ~w6137;
assign w6149 = ~w6147 & w6148;
assign w6150 = ~w6142 & ~w6144;
assign w6151 = ~w6149 & ~w6150;
assign w6152 = w6148 & w6147;
assign w6153 = ~w6147 & ~w6148;
assign w6154 = ~w6152 & ~w6153;
assign w6155 = ~w6151 & ~w6154;
assign w6156 = ~w6140 & ~w6155;
assign w6157 = ~A_115 & A_116;
assign w6158 = A_115 & ~A_116;
assign w6159 = A_117 & ~w6158;
assign w6160 = ~w6157 & w6159;
assign w6161 = ~w6157 & ~w6158;
assign w6162 = ~A_117 & ~w6161;
assign w6163 = ~w6160 & ~w6162;
assign w6164 = ~A_118 & A_119;
assign w6165 = A_118 & ~A_119;
assign w6166 = A_120 & ~w6165;
assign w6167 = ~w6164 & w6166;
assign w6168 = ~w6164 & ~w6165;
assign w6169 = ~A_120 & ~w6168;
assign w6170 = ~w6167 & ~w6169;
assign w6171 = ~w6163 & w6170;
assign w6172 = w6163 & ~w6170;
assign w6173 = ~w6171 & ~w6172;
assign w6174 = A_118 & A_119;
assign w6175 = (~w6174 & w6168) | (~w6174 & w12774) | (w6168 & w12774);
assign w6176 = A_115 & A_116;
assign w6177 = (~w6176 & w6161) | (~w6176 & w12775) | (w6161 & w12775);
assign w6178 = ~w6175 & w6177;
assign w6179 = w6175 & ~w6177;
assign w6180 = ~w6178 & ~w6179;
assign w6181 = ~w6163 & ~w6170;
assign w6182 = ~w6180 & w6181;
assign w6183 = ~w6175 & ~w6177;
assign w6184 = ~w6182 & ~w6183;
assign w6185 = w6181 & w6180;
assign w6186 = ~w6180 & ~w6181;
assign w6187 = ~w6185 & ~w6186;
assign w6188 = ~w6184 & ~w6187;
assign w6189 = ~w6173 & ~w6188;
assign w6190 = ~w6156 & w6189;
assign w6191 = w6156 & ~w6189;
assign w6192 = ~w6190 & ~w6191;
assign w6193 = ~A_109 & A_110;
assign w6194 = A_109 & ~A_110;
assign w6195 = A_111 & ~w6194;
assign w6196 = ~w6193 & w6195;
assign w6197 = ~w6193 & ~w6194;
assign w6198 = ~A_111 & ~w6197;
assign w6199 = ~w6196 & ~w6198;
assign w6200 = ~A_112 & A_113;
assign w6201 = A_112 & ~A_113;
assign w6202 = A_114 & ~w6201;
assign w6203 = ~w6200 & w6202;
assign w6204 = ~w6200 & ~w6201;
assign w6205 = ~A_114 & ~w6204;
assign w6206 = ~w6203 & ~w6205;
assign w6207 = ~w6199 & w6206;
assign w6208 = w6199 & ~w6206;
assign w6209 = ~w6207 & ~w6208;
assign w6210 = A_112 & A_113;
assign w6211 = (~w6210 & w6204) | (~w6210 & w12776) | (w6204 & w12776);
assign w6212 = A_109 & A_110;
assign w6213 = (~w6212 & w6197) | (~w6212 & w12777) | (w6197 & w12777);
assign w6214 = ~w6211 & w6213;
assign w6215 = w6211 & ~w6213;
assign w6216 = ~w6214 & ~w6215;
assign w6217 = ~w6199 & ~w6206;
assign w6218 = ~w6216 & w6217;
assign w6219 = ~w6211 & ~w6213;
assign w6220 = ~w6218 & ~w6219;
assign w6221 = w6217 & w6216;
assign w6222 = ~w6216 & ~w6217;
assign w6223 = ~w6221 & ~w6222;
assign w6224 = ~w6220 & ~w6223;
assign w6225 = ~w6209 & ~w6224;
assign w6226 = ~A_103 & A_104;
assign w6227 = A_103 & ~A_104;
assign w6228 = A_105 & ~w6227;
assign w6229 = ~w6226 & w6228;
assign w6230 = ~w6226 & ~w6227;
assign w6231 = ~A_105 & ~w6230;
assign w6232 = ~w6229 & ~w6231;
assign w6233 = ~A_106 & A_107;
assign w6234 = A_106 & ~A_107;
assign w6235 = A_108 & ~w6234;
assign w6236 = ~w6233 & w6235;
assign w6237 = ~w6233 & ~w6234;
assign w6238 = ~A_108 & ~w6237;
assign w6239 = ~w6236 & ~w6238;
assign w6240 = ~w6232 & w6239;
assign w6241 = w6232 & ~w6239;
assign w6242 = ~w6240 & ~w6241;
assign w6243 = A_106 & A_107;
assign w6244 = (~w6243 & w6237) | (~w6243 & w12778) | (w6237 & w12778);
assign w6245 = A_103 & A_104;
assign w6246 = (~w6245 & w6230) | (~w6245 & w12779) | (w6230 & w12779);
assign w6247 = ~w6244 & w6246;
assign w6248 = w6244 & ~w6246;
assign w6249 = ~w6247 & ~w6248;
assign w6250 = ~w6232 & ~w6239;
assign w6251 = ~w6249 & w6250;
assign w6252 = ~w6244 & ~w6246;
assign w6253 = ~w6251 & ~w6252;
assign w6254 = w6250 & w6249;
assign w6255 = ~w6249 & ~w6250;
assign w6256 = ~w6254 & ~w6255;
assign w6257 = ~w6253 & ~w6256;
assign w6258 = ~w6242 & ~w6257;
assign w6259 = ~w6225 & w6258;
assign w6260 = w6225 & ~w6258;
assign w6261 = ~w6259 & ~w6260;
assign w6262 = ~w6192 & w6261;
assign w6263 = w6192 & ~w6261;
assign w6264 = ~w6262 & ~w6263;
assign w6265 = ~A_97 & A_98;
assign w6266 = A_97 & ~A_98;
assign w6267 = A_99 & ~w6266;
assign w6268 = ~w6265 & w6267;
assign w6269 = ~w6265 & ~w6266;
assign w6270 = ~A_99 & ~w6269;
assign w6271 = ~w6268 & ~w6270;
assign w6272 = ~A_100 & A_101;
assign w6273 = A_100 & ~A_101;
assign w6274 = A_102 & ~w6273;
assign w6275 = ~w6272 & w6274;
assign w6276 = ~w6272 & ~w6273;
assign w6277 = ~A_102 & ~w6276;
assign w6278 = ~w6275 & ~w6277;
assign w6279 = ~w6271 & w6278;
assign w6280 = w6271 & ~w6278;
assign w6281 = ~w6279 & ~w6280;
assign w6282 = A_100 & A_101;
assign w6283 = (~w6282 & w6276) | (~w6282 & w12780) | (w6276 & w12780);
assign w6284 = A_97 & A_98;
assign w6285 = (~w6284 & w6269) | (~w6284 & w12781) | (w6269 & w12781);
assign w6286 = ~w6283 & w6285;
assign w6287 = w6283 & ~w6285;
assign w6288 = ~w6286 & ~w6287;
assign w6289 = ~w6271 & ~w6278;
assign w6290 = ~w6288 & w6289;
assign w6291 = ~w6283 & ~w6285;
assign w6292 = ~w6290 & ~w6291;
assign w6293 = w6289 & w6288;
assign w6294 = ~w6288 & ~w6289;
assign w6295 = ~w6293 & ~w6294;
assign w6296 = ~w6292 & ~w6295;
assign w6297 = ~w6281 & ~w6296;
assign w6298 = ~A_91 & A_92;
assign w6299 = A_91 & ~A_92;
assign w6300 = A_93 & ~w6299;
assign w6301 = ~w6298 & w6300;
assign w6302 = ~w6298 & ~w6299;
assign w6303 = ~A_93 & ~w6302;
assign w6304 = ~w6301 & ~w6303;
assign w6305 = ~A_94 & A_95;
assign w6306 = A_94 & ~A_95;
assign w6307 = A_96 & ~w6306;
assign w6308 = ~w6305 & w6307;
assign w6309 = ~w6305 & ~w6306;
assign w6310 = ~A_96 & ~w6309;
assign w6311 = ~w6308 & ~w6310;
assign w6312 = ~w6304 & w6311;
assign w6313 = w6304 & ~w6311;
assign w6314 = ~w6312 & ~w6313;
assign w6315 = A_94 & A_95;
assign w6316 = (~w6315 & w6309) | (~w6315 & w12782) | (w6309 & w12782);
assign w6317 = A_91 & A_92;
assign w6318 = (~w6317 & w6302) | (~w6317 & w12783) | (w6302 & w12783);
assign w6319 = ~w6316 & w6318;
assign w6320 = w6316 & ~w6318;
assign w6321 = ~w6319 & ~w6320;
assign w6322 = ~w6304 & ~w6311;
assign w6323 = ~w6321 & w6322;
assign w6324 = ~w6316 & ~w6318;
assign w6325 = ~w6323 & ~w6324;
assign w6326 = w6322 & w6321;
assign w6327 = ~w6321 & ~w6322;
assign w6328 = ~w6326 & ~w6327;
assign w6329 = ~w6325 & ~w6328;
assign w6330 = ~w6314 & ~w6329;
assign w6331 = ~w6297 & w6330;
assign w6332 = w6297 & ~w6330;
assign w6333 = ~w6331 & ~w6332;
assign w6334 = ~A_85 & A_86;
assign w6335 = A_85 & ~A_86;
assign w6336 = A_87 & ~w6335;
assign w6337 = ~w6334 & w6336;
assign w6338 = ~w6334 & ~w6335;
assign w6339 = ~A_87 & ~w6338;
assign w6340 = ~w6337 & ~w6339;
assign w6341 = ~A_88 & A_89;
assign w6342 = A_88 & ~A_89;
assign w6343 = A_90 & ~w6342;
assign w6344 = ~w6341 & w6343;
assign w6345 = ~w6341 & ~w6342;
assign w6346 = ~A_90 & ~w6345;
assign w6347 = ~w6344 & ~w6346;
assign w6348 = ~w6340 & w6347;
assign w6349 = w6340 & ~w6347;
assign w6350 = ~w6348 & ~w6349;
assign w6351 = A_88 & A_89;
assign w6352 = (~w6351 & w6345) | (~w6351 & w12784) | (w6345 & w12784);
assign w6353 = A_85 & A_86;
assign w6354 = (~w6353 & w6338) | (~w6353 & w12785) | (w6338 & w12785);
assign w6355 = ~w6352 & w6354;
assign w6356 = w6352 & ~w6354;
assign w6357 = ~w6355 & ~w6356;
assign w6358 = ~w6340 & ~w6347;
assign w6359 = ~w6357 & w6358;
assign w6360 = ~w6352 & ~w6354;
assign w6361 = ~w6359 & ~w6360;
assign w6362 = w6358 & w6357;
assign w6363 = ~w6357 & ~w6358;
assign w6364 = ~w6362 & ~w6363;
assign w6365 = ~w6361 & ~w6364;
assign w6366 = ~w6350 & ~w6365;
assign w6367 = ~A_79 & A_80;
assign w6368 = A_79 & ~A_80;
assign w6369 = A_81 & ~w6368;
assign w6370 = ~w6367 & w6369;
assign w6371 = ~w6367 & ~w6368;
assign w6372 = ~A_81 & ~w6371;
assign w6373 = ~w6370 & ~w6372;
assign w6374 = ~A_82 & A_83;
assign w6375 = A_82 & ~A_83;
assign w6376 = A_84 & ~w6375;
assign w6377 = ~w6374 & w6376;
assign w6378 = ~w6374 & ~w6375;
assign w6379 = ~A_84 & ~w6378;
assign w6380 = ~w6377 & ~w6379;
assign w6381 = ~w6373 & w6380;
assign w6382 = w6373 & ~w6380;
assign w6383 = ~w6381 & ~w6382;
assign w6384 = A_82 & A_83;
assign w6385 = (~w6384 & w6378) | (~w6384 & w12786) | (w6378 & w12786);
assign w6386 = A_79 & A_80;
assign w6387 = (~w6386 & w6371) | (~w6386 & w12787) | (w6371 & w12787);
assign w6388 = ~w6385 & w6387;
assign w6389 = w6385 & ~w6387;
assign w6390 = ~w6388 & ~w6389;
assign w6391 = ~w6373 & ~w6380;
assign w6392 = ~w6390 & w6391;
assign w6393 = ~w6385 & ~w6387;
assign w6394 = ~w6392 & ~w6393;
assign w6395 = w6391 & w6390;
assign w6396 = ~w6390 & ~w6391;
assign w6397 = ~w6395 & ~w6396;
assign w6398 = ~w6394 & ~w6397;
assign w6399 = ~w6383 & ~w6398;
assign w6400 = ~w6366 & w6399;
assign w6401 = w6366 & ~w6399;
assign w6402 = ~w6400 & ~w6401;
assign w6403 = ~w6333 & w6402;
assign w6404 = w6333 & ~w6402;
assign w6405 = ~w6403 & ~w6404;
assign w6406 = ~w6264 & w6405;
assign w6407 = w6264 & ~w6405;
assign w6408 = ~w6406 & ~w6407;
assign w6409 = ~w6123 & w6408;
assign w6410 = w6123 & ~w6408;
assign w6411 = ~w6409 & ~w6410;
assign w6412 = ~w5838 & ~w6411;
assign w6413 = (w6412 & w5834) | (w6412 & w13873) | (w5834 & w13873);
assign w6414 = ~w5830 & w6413;
assign w6415 = ~w5830 & ~w5835;
assign w6416 = ~w6412 & ~w6415;
assign w6417 = ~w6029 & ~w6040;
assign w6418 = ~w6043 & ~w6417;
assign w6419 = ~w5996 & ~w6029;
assign w6420 = ~w6011 & w6419;
assign w6421 = ~w6044 & w6420;
assign w6422 = ~w5996 & ~w6007;
assign w6423 = ~w6010 & ~w6422;
assign w6424 = ~w6421 & ~w6423;
assign w6425 = ~w6010 & w6419;
assign w6426 = ~w6011 & w6425;
assign w6427 = ~w6044 & ~w6422;
assign w6428 = w6426 & w6427;
assign w6429 = (w6418 & w6424) | (w6418 & w12998) | (w6424 & w12998);
assign w6430 = ~w6421 & w6423;
assign w6431 = w6421 & ~w6423;
assign w6432 = ~w6430 & ~w6431;
assign w6433 = ~w6418 & ~w6432;
assign w6434 = ~w6048 & ~w6117;
assign w6435 = ~w6433 & w13382;
assign w6436 = (~w6434 & w6433) | (~w6434 & w13383) | (w6433 & w13383);
assign w6437 = ~w6435 & ~w6436;
assign w6438 = ~w6098 & ~w6109;
assign w6439 = ~w6112 & ~w6438;
assign w6440 = ~w6065 & ~w6098;
assign w6441 = ~w6080 & w6440;
assign w6442 = ~w6113 & w6441;
assign w6443 = ~w6065 & ~w6076;
assign w6444 = ~w6079 & ~w6443;
assign w6445 = ~w6442 & w6444;
assign w6446 = w6442 & ~w6444;
assign w6447 = ~w6445 & ~w6446;
assign w6448 = ~w6439 & ~w6447;
assign w6449 = ~w6442 & ~w6444;
assign w6450 = ~w6079 & w6440;
assign w6451 = ~w6080 & w6450;
assign w6452 = ~w6113 & ~w6443;
assign w6453 = w6451 & w6452;
assign w6454 = (w6439 & w6449) | (w6439 & w13384) | (w6449 & w13384);
assign w6455 = ~w6448 & ~w6454;
assign w6456 = ~w6437 & w6455;
assign w6457 = ~w6433 & w12999;
assign w6458 = (w6434 & w6433) | (w6434 & w13385) | (w6433 & w13385);
assign w6459 = ~w6457 & ~w6458;
assign w6460 = ~w6455 & ~w6459;
assign w6461 = ~w6456 & ~w6460;
assign w6462 = ~w5957 & ~w5968;
assign w6463 = ~w5971 & ~w6462;
assign w6464 = ~w5924 & ~w5957;
assign w6465 = ~w5939 & w6464;
assign w6466 = ~w5972 & w6465;
assign w6467 = ~w5924 & ~w5935;
assign w6468 = ~w5938 & ~w6467;
assign w6469 = ~w6466 & w6468;
assign w6470 = w6466 & ~w6468;
assign w6471 = ~w6469 & ~w6470;
assign w6472 = ~w6463 & ~w6471;
assign w6473 = ~w6466 & ~w6468;
assign w6474 = ~w5938 & w6464;
assign w6475 = ~w5939 & w6474;
assign w6476 = ~w5972 & ~w6467;
assign w6477 = w6475 & w6476;
assign w6478 = (w6463 & w6473) | (w6463 & w13386) | (w6473 & w13386);
assign w6479 = ~w6472 & ~w6478;
assign w6480 = ~w5888 & ~w5899;
assign w6481 = ~w5902 & ~w6480;
assign w6482 = ~w5855 & ~w5888;
assign w6483 = ~w5870 & w6482;
assign w6484 = ~w5903 & w6483;
assign w6485 = ~w5855 & ~w5866;
assign w6486 = ~w5869 & ~w6485;
assign w6487 = ~w6484 & ~w6486;
assign w6488 = ~w5869 & w6482;
assign w6489 = ~w5870 & w6488;
assign w6490 = ~w5903 & ~w6485;
assign w6491 = w6489 & w6490;
assign w6492 = (w6481 & w6487) | (w6481 & w13000) | (w6487 & w13000);
assign w6493 = ~w6484 & w6486;
assign w6494 = w6484 & ~w6486;
assign w6495 = ~w6493 & ~w6494;
assign w6496 = ~w6481 & ~w6495;
assign w6497 = ~w5907 & ~w5976;
assign w6498 = ~w6496 & w13001;
assign w6499 = (w6497 & w6496) | (w6497 & w13002) | (w6496 & w13002);
assign w6500 = ~w6498 & ~w6499;
assign w6501 = ~w6479 & ~w6500;
assign w6502 = ~w6496 & w13003;
assign w6503 = (~w6497 & w6496) | (~w6497 & w13387) | (w6496 & w13387);
assign w6504 = (w6479 & w6503) | (w6479 & w13004) | (w6503 & w13004);
assign w6505 = ~w5979 & ~w6120;
assign w6506 = ~w6505 & ~w6504;
assign w6507 = ~w6501 & w6506;
assign w6508 = ~w6501 & ~w6504;
assign w6509 = w6505 & ~w6508;
assign w6510 = (~w6461 & w6509) | (~w6461 & w13874) | (w6509 & w13874);
assign w6511 = w6505 & ~w6504;
assign w6512 = ~w6501 & w6511;
assign w6513 = ~w6505 & ~w6508;
assign w6514 = (w6461 & w6513) | (w6461 & w13388) | (w6513 & w13388);
assign w6515 = ~w6123 & ~w6408;
assign w6516 = ~w6514 & w6515;
assign w6517 = ~w6510 & w6516;
assign w6518 = ~w6510 & ~w6514;
assign w6519 = ~w6515 & ~w6518;
assign w6520 = ~w6517 & ~w6519;
assign w6521 = ~w6242 & ~w6253;
assign w6522 = ~w6256 & ~w6521;
assign w6523 = ~w6209 & ~w6242;
assign w6524 = ~w6224 & w6523;
assign w6525 = ~w6257 & w6524;
assign w6526 = ~w6209 & ~w6220;
assign w6527 = ~w6223 & ~w6526;
assign w6528 = ~w6525 & w6527;
assign w6529 = w6525 & ~w6527;
assign w6530 = ~w6528 & ~w6529;
assign w6531 = ~w6522 & ~w6530;
assign w6532 = ~w6525 & ~w6527;
assign w6533 = ~w6223 & w6523;
assign w6534 = ~w6224 & w6533;
assign w6535 = ~w6257 & ~w6526;
assign w6536 = w6534 & w6535;
assign w6537 = (w6522 & w6532) | (w6522 & w13389) | (w6532 & w13389);
assign w6538 = ~w6531 & ~w6537;
assign w6539 = ~w6173 & ~w6184;
assign w6540 = ~w6187 & ~w6539;
assign w6541 = ~w6140 & ~w6173;
assign w6542 = ~w6155 & w6541;
assign w6543 = ~w6188 & w6542;
assign w6544 = ~w6140 & ~w6151;
assign w6545 = ~w6154 & ~w6544;
assign w6546 = ~w6543 & ~w6545;
assign w6547 = ~w6154 & w6541;
assign w6548 = ~w6155 & w6547;
assign w6549 = ~w6188 & ~w6544;
assign w6550 = w6548 & w6549;
assign w6551 = (w6540 & w6546) | (w6540 & w13005) | (w6546 & w13005);
assign w6552 = ~w6543 & w6545;
assign w6553 = w6543 & ~w6545;
assign w6554 = ~w6552 & ~w6553;
assign w6555 = ~w6540 & ~w6554;
assign w6556 = ~w6192 & ~w6261;
assign w6557 = ~w6555 & w13006;
assign w6558 = (w6556 & w6555) | (w6556 & w13007) | (w6555 & w13007);
assign w6559 = ~w6557 & ~w6558;
assign w6560 = ~w6538 & ~w6559;
assign w6561 = ~w6555 & w13008;
assign w6562 = (~w6556 & w6555) | (~w6556 & w13390) | (w6555 & w13390);
assign w6563 = (w6538 & w6562) | (w6538 & w13009) | (w6562 & w13009);
assign w6564 = ~w6264 & ~w6405;
assign w6565 = w6564 & ~w6563;
assign w6566 = ~w6560 & w6565;
assign w6567 = ~w6560 & ~w6563;
assign w6568 = ~w6564 & ~w6567;
assign w6569 = ~w6314 & ~w6325;
assign w6570 = ~w6328 & ~w6569;
assign w6571 = ~w6281 & ~w6314;
assign w6572 = ~w6296 & w6571;
assign w6573 = ~w6329 & w6572;
assign w6574 = ~w6281 & ~w6292;
assign w6575 = ~w6295 & ~w6574;
assign w6576 = ~w6573 & ~w6575;
assign w6577 = ~w6295 & w6571;
assign w6578 = ~w6296 & w6577;
assign w6579 = ~w6329 & ~w6574;
assign w6580 = w6578 & w6579;
assign w6581 = (w6570 & w6576) | (w6570 & w13010) | (w6576 & w13010);
assign w6582 = ~w6573 & w6575;
assign w6583 = w6573 & ~w6575;
assign w6584 = ~w6582 & ~w6583;
assign w6585 = ~w6570 & ~w6584;
assign w6586 = ~w6333 & ~w6402;
assign w6587 = ~w6585 & w13391;
assign w6588 = (~w6586 & w6585) | (~w6586 & w13392) | (w6585 & w13392);
assign w6589 = ~w6587 & ~w6588;
assign w6590 = ~w6383 & ~w6394;
assign w6591 = ~w6397 & ~w6590;
assign w6592 = ~w6350 & ~w6383;
assign w6593 = ~w6365 & w6592;
assign w6594 = ~w6398 & w6593;
assign w6595 = ~w6350 & ~w6361;
assign w6596 = ~w6364 & ~w6595;
assign w6597 = ~w6594 & w6596;
assign w6598 = w6594 & ~w6596;
assign w6599 = ~w6597 & ~w6598;
assign w6600 = ~w6591 & ~w6599;
assign w6601 = ~w6594 & ~w6596;
assign w6602 = ~w6364 & w6592;
assign w6603 = ~w6365 & w6602;
assign w6604 = ~w6398 & ~w6595;
assign w6605 = w6603 & w6604;
assign w6606 = (w6591 & w6601) | (w6591 & w13393) | (w6601 & w13393);
assign w6607 = ~w6600 & ~w6606;
assign w6608 = ~w6589 & w6607;
assign w6609 = ~w6585 & w13011;
assign w6610 = (w6586 & w6585) | (w6586 & w13394) | (w6585 & w13394);
assign w6611 = ~w6609 & ~w6610;
assign w6612 = ~w6607 & ~w6611;
assign w6613 = ~w6608 & ~w6612;
assign w6614 = (w6613 & w6568) | (w6613 & w13875) | (w6568 & w13875);
assign w6615 = ~w6564 & ~w6563;
assign w6616 = ~w6560 & w6615;
assign w6617 = w6564 & ~w6567;
assign w6618 = (~w6613 & w6617) | (~w6613 & w13876) | (w6617 & w13876);
assign w6619 = ~w6614 & ~w6618;
assign w6620 = ~w6520 & w6619;
assign w6621 = ~w6514 & ~w6515;
assign w6622 = ~w6510 & w6621;
assign w6623 = w6515 & ~w6518;
assign w6624 = ~w6622 & ~w6623;
assign w6625 = ~w6619 & ~w6624;
assign w6626 = ~w6620 & ~w6625;
assign w6627 = (w6626 & w6416) | (w6626 & w13877) | (w6416 & w13877);
assign w6628 = (~w6412 & w5834) | (~w6412 & w14063) | (w5834 & w14063);
assign w6629 = ~w5830 & w6628;
assign w6630 = w6412 & ~w6415;
assign w6631 = (~w6626 & w6630) | (~w6626 & w14064) | (w6630 & w14064);
assign w6632 = ~w6627 & ~w6631;
assign w6633 = A_334 & A_335;
assign w6634 = A_334 & ~A_335;
assign w6635 = ~A_334 & A_335;
assign w6636 = ~w6634 & ~w6635;
assign w6637 = (~w6633 & w6636) | (~w6633 & w12788) | (w6636 & w12788);
assign w6638 = A_331 & A_332;
assign w6639 = A_331 & ~A_332;
assign w6640 = ~A_331 & A_332;
assign w6641 = ~w6639 & ~w6640;
assign w6642 = (~w6638 & w6641) | (~w6638 & w12789) | (w6641 & w12789);
assign w6643 = w6637 & ~w6642;
assign w6644 = ~w6637 & w6642;
assign w6645 = A_333 & ~w6639;
assign w6646 = ~w6640 & w6645;
assign w6647 = ~A_333 & ~w6641;
assign w6648 = ~w6646 & ~w6647;
assign w6649 = A_336 & ~w6634;
assign w6650 = ~w6635 & w6649;
assign w6651 = ~A_336 & ~w6636;
assign w6652 = ~w6650 & ~w6651;
assign w6653 = ~w6648 & ~w6652;
assign w6654 = w6653 & w6655;
assign w6655 = ~w6643 & ~w6644;
assign w6656 = ~w6653 & ~w6655;
assign w6657 = ~w6654 & ~w6656;
assign w6658 = ~w6648 & w6652;
assign w6659 = w6648 & ~w6652;
assign w6660 = ~w6658 & ~w6659;
assign w6661 = w6653 & ~w6655;
assign w6662 = ~w6637 & ~w6642;
assign w6663 = ~w6661 & ~w6662;
assign w6664 = ~w6660 & ~w6663;
assign w6665 = ~w6657 & ~w6664;
assign w6666 = ~w6657 & ~w6663;
assign w6667 = A_340 & A_341;
assign w6668 = A_340 & ~A_341;
assign w6669 = ~A_340 & A_341;
assign w6670 = ~w6668 & ~w6669;
assign w6671 = (~w6667 & w6670) | (~w6667 & w12790) | (w6670 & w12790);
assign w6672 = A_337 & A_338;
assign w6673 = A_337 & ~A_338;
assign w6674 = ~A_337 & A_338;
assign w6675 = ~w6673 & ~w6674;
assign w6676 = (~w6672 & w6675) | (~w6672 & w12791) | (w6675 & w12791);
assign w6677 = ~w6671 & w6676;
assign w6678 = w6671 & ~w6676;
assign w6679 = ~w6677 & ~w6678;
assign w6680 = A_339 & ~w6673;
assign w6681 = ~w6674 & w6680;
assign w6682 = ~A_339 & ~w6675;
assign w6683 = ~w6681 & ~w6682;
assign w6684 = A_342 & ~w6668;
assign w6685 = ~w6669 & w6684;
assign w6686 = ~A_342 & ~w6670;
assign w6687 = ~w6685 & ~w6686;
assign w6688 = ~w6683 & ~w6687;
assign w6689 = ~w6679 & w6688;
assign w6690 = ~w6671 & ~w6676;
assign w6691 = ~w6689 & ~w6690;
assign w6692 = w6688 & w6679;
assign w6693 = ~w6679 & ~w6688;
assign w6694 = ~w6692 & ~w6693;
assign w6695 = ~w6691 & ~w6694;
assign w6696 = ~w6683 & w6687;
assign w6697 = w6683 & ~w6687;
assign w6698 = ~w6696 & ~w6697;
assign w6699 = ~w6660 & ~w6698;
assign w6700 = ~w6695 & w6699;
assign w6701 = ~w6666 & w6700;
assign w6702 = ~w6691 & ~w6698;
assign w6703 = ~w6694 & ~w6702;
assign w6704 = ~w6701 & ~w6703;
assign w6705 = ~w6694 & w6699;
assign w6706 = ~w6695 & w6705;
assign w6707 = ~w6666 & ~w6702;
assign w6708 = w6706 & w6707;
assign w6709 = (w6665 & w6704) | (w6665 & w13012) | (w6704 & w13012);
assign w6710 = ~w6701 & w6703;
assign w6711 = w6701 & ~w6703;
assign w6712 = ~w6710 & ~w6711;
assign w6713 = ~w6665 & ~w6712;
assign w6714 = ~w6695 & ~w6698;
assign w6715 = ~w6660 & ~w6666;
assign w6716 = ~w6714 & w6715;
assign w6717 = w6714 & ~w6715;
assign w6718 = ~w6716 & ~w6717;
assign w6719 = ~A_325 & A_326;
assign w6720 = A_325 & ~A_326;
assign w6721 = A_327 & ~w6720;
assign w6722 = ~w6719 & w6721;
assign w6723 = ~w6719 & ~w6720;
assign w6724 = ~A_327 & ~w6723;
assign w6725 = ~w6722 & ~w6724;
assign w6726 = ~A_328 & A_329;
assign w6727 = A_328 & ~A_329;
assign w6728 = A_330 & ~w6727;
assign w6729 = ~w6726 & w6728;
assign w6730 = ~w6726 & ~w6727;
assign w6731 = ~A_330 & ~w6730;
assign w6732 = ~w6729 & ~w6731;
assign w6733 = ~w6725 & w6732;
assign w6734 = w6725 & ~w6732;
assign w6735 = ~w6733 & ~w6734;
assign w6736 = A_328 & A_329;
assign w6737 = (~w6736 & w6730) | (~w6736 & w12792) | (w6730 & w12792);
assign w6738 = A_325 & A_326;
assign w6739 = (~w6738 & w6723) | (~w6738 & w12793) | (w6723 & w12793);
assign w6740 = ~w6737 & w6739;
assign w6741 = w6737 & ~w6739;
assign w6742 = ~w6740 & ~w6741;
assign w6743 = ~w6725 & ~w6732;
assign w6744 = ~w6742 & w6743;
assign w6745 = ~w6737 & ~w6739;
assign w6746 = ~w6744 & ~w6745;
assign w6747 = w6743 & w6742;
assign w6748 = ~w6742 & ~w6743;
assign w6749 = ~w6747 & ~w6748;
assign w6750 = ~w6746 & ~w6749;
assign w6751 = ~w6735 & ~w6750;
assign w6752 = ~A_319 & A_320;
assign w6753 = A_319 & ~A_320;
assign w6754 = A_321 & ~w6753;
assign w6755 = ~w6752 & w6754;
assign w6756 = ~w6752 & ~w6753;
assign w6757 = ~A_321 & ~w6756;
assign w6758 = ~w6755 & ~w6757;
assign w6759 = ~A_322 & A_323;
assign w6760 = A_322 & ~A_323;
assign w6761 = A_324 & ~w6760;
assign w6762 = ~w6759 & w6761;
assign w6763 = ~w6759 & ~w6760;
assign w6764 = ~A_324 & ~w6763;
assign w6765 = ~w6762 & ~w6764;
assign w6766 = ~w6758 & w6765;
assign w6767 = w6758 & ~w6765;
assign w6768 = ~w6766 & ~w6767;
assign w6769 = A_322 & A_323;
assign w6770 = (~w6769 & w6763) | (~w6769 & w12794) | (w6763 & w12794);
assign w6771 = A_319 & A_320;
assign w6772 = (~w6771 & w6756) | (~w6771 & w12795) | (w6756 & w12795);
assign w6773 = ~w6770 & w6772;
assign w6774 = w6770 & ~w6772;
assign w6775 = ~w6773 & ~w6774;
assign w6776 = ~w6758 & ~w6765;
assign w6777 = ~w6775 & w6776;
assign w6778 = ~w6770 & ~w6772;
assign w6779 = ~w6777 & ~w6778;
assign w6780 = w6776 & w6775;
assign w6781 = ~w6775 & ~w6776;
assign w6782 = ~w6780 & ~w6781;
assign w6783 = ~w6779 & ~w6782;
assign w6784 = ~w6768 & ~w6783;
assign w6785 = ~w6751 & w6784;
assign w6786 = w6751 & ~w6784;
assign w6787 = ~w6785 & ~w6786;
assign w6788 = ~w6718 & ~w6787;
assign w6789 = ~w6713 & w13395;
assign w6790 = (~w6788 & w6713) | (~w6788 & w13396) | (w6713 & w13396);
assign w6791 = ~w6789 & ~w6790;
assign w6792 = ~w6768 & ~w6779;
assign w6793 = ~w6782 & ~w6792;
assign w6794 = ~w6735 & ~w6768;
assign w6795 = ~w6750 & w6794;
assign w6796 = ~w6783 & w6795;
assign w6797 = ~w6735 & ~w6746;
assign w6798 = ~w6749 & ~w6797;
assign w6799 = ~w6796 & w6798;
assign w6800 = w6796 & ~w6798;
assign w6801 = ~w6799 & ~w6800;
assign w6802 = ~w6793 & ~w6801;
assign w6803 = ~w6796 & ~w6798;
assign w6804 = ~w6749 & w6794;
assign w6805 = ~w6750 & w6804;
assign w6806 = ~w6783 & ~w6797;
assign w6807 = w6805 & w6806;
assign w6808 = (w6793 & w6803) | (w6793 & w13397) | (w6803 & w13397);
assign w6809 = ~w6802 & ~w6808;
assign w6810 = ~w6791 & w6809;
assign w6811 = ~w6713 & w13013;
assign w6812 = (w6788 & w6713) | (w6788 & w13398) | (w6713 & w13398);
assign w6813 = ~w6811 & ~w6812;
assign w6814 = ~w6809 & ~w6813;
assign w6815 = ~w6810 & ~w6814;
assign w6816 = A_346 & A_347;
assign w6817 = A_346 & ~A_347;
assign w6818 = ~A_346 & A_347;
assign w6819 = ~w6817 & ~w6818;
assign w6820 = (~w6816 & w6819) | (~w6816 & w12796) | (w6819 & w12796);
assign w6821 = A_343 & A_344;
assign w6822 = A_343 & ~A_344;
assign w6823 = ~A_343 & A_344;
assign w6824 = ~w6822 & ~w6823;
assign w6825 = (~w6821 & w6824) | (~w6821 & w12797) | (w6824 & w12797);
assign w6826 = w6820 & ~w6825;
assign w6827 = ~w6820 & w6825;
assign w6828 = A_345 & ~w6822;
assign w6829 = ~w6823 & w6828;
assign w6830 = ~A_345 & ~w6824;
assign w6831 = ~w6829 & ~w6830;
assign w6832 = A_348 & ~w6817;
assign w6833 = ~w6818 & w6832;
assign w6834 = ~A_348 & ~w6819;
assign w6835 = ~w6833 & ~w6834;
assign w6836 = ~w6831 & ~w6835;
assign w6837 = w6836 & w6838;
assign w6838 = ~w6826 & ~w6827;
assign w6839 = ~w6836 & ~w6838;
assign w6840 = ~w6837 & ~w6839;
assign w6841 = ~w6831 & w6835;
assign w6842 = w6831 & ~w6835;
assign w6843 = ~w6841 & ~w6842;
assign w6844 = w6836 & ~w6838;
assign w6845 = ~w6820 & ~w6825;
assign w6846 = ~w6844 & ~w6845;
assign w6847 = ~w6843 & ~w6846;
assign w6848 = ~w6840 & ~w6847;
assign w6849 = ~w6840 & ~w6846;
assign w6850 = A_352 & A_353;
assign w6851 = A_352 & ~A_353;
assign w6852 = ~A_352 & A_353;
assign w6853 = ~w6851 & ~w6852;
assign w6854 = (~w6850 & w6853) | (~w6850 & w12798) | (w6853 & w12798);
assign w6855 = A_349 & A_350;
assign w6856 = A_349 & ~A_350;
assign w6857 = ~A_349 & A_350;
assign w6858 = ~w6856 & ~w6857;
assign w6859 = (~w6855 & w6858) | (~w6855 & w12799) | (w6858 & w12799);
assign w6860 = ~w6854 & w6859;
assign w6861 = w6854 & ~w6859;
assign w6862 = ~w6860 & ~w6861;
assign w6863 = A_351 & ~w6856;
assign w6864 = ~w6857 & w6863;
assign w6865 = ~A_351 & ~w6858;
assign w6866 = ~w6864 & ~w6865;
assign w6867 = A_354 & ~w6851;
assign w6868 = ~w6852 & w6867;
assign w6869 = ~A_354 & ~w6853;
assign w6870 = ~w6868 & ~w6869;
assign w6871 = ~w6866 & ~w6870;
assign w6872 = ~w6862 & w6871;
assign w6873 = ~w6854 & ~w6859;
assign w6874 = ~w6872 & ~w6873;
assign w6875 = w6871 & w6862;
assign w6876 = ~w6862 & ~w6871;
assign w6877 = ~w6875 & ~w6876;
assign w6878 = ~w6874 & ~w6877;
assign w6879 = ~w6866 & w6870;
assign w6880 = w6866 & ~w6870;
assign w6881 = ~w6879 & ~w6880;
assign w6882 = ~w6843 & ~w6881;
assign w6883 = ~w6878 & w6882;
assign w6884 = ~w6849 & w6883;
assign w6885 = ~w6874 & ~w6881;
assign w6886 = ~w6877 & ~w6885;
assign w6887 = ~w6884 & w6886;
assign w6888 = w6884 & ~w6886;
assign w6889 = ~w6887 & ~w6888;
assign w6890 = ~w6848 & ~w6889;
assign w6891 = ~w6884 & ~w6886;
assign w6892 = ~w6877 & w6882;
assign w6893 = ~w6878 & w6892;
assign w6894 = ~w6849 & ~w6885;
assign w6895 = w6893 & w6894;
assign w6896 = (w6848 & w6891) | (w6848 & w13399) | (w6891 & w13399);
assign w6897 = ~w6890 & ~w6896;
assign w6898 = A_358 & A_359;
assign w6899 = A_358 & ~A_359;
assign w6900 = ~A_358 & A_359;
assign w6901 = ~w6899 & ~w6900;
assign w6902 = (~w6898 & w6901) | (~w6898 & w12800) | (w6901 & w12800);
assign w6903 = A_355 & A_356;
assign w6904 = A_355 & ~A_356;
assign w6905 = ~A_355 & A_356;
assign w6906 = ~w6904 & ~w6905;
assign w6907 = (~w6903 & w6906) | (~w6903 & w12801) | (w6906 & w12801);
assign w6908 = w6902 & ~w6907;
assign w6909 = ~w6902 & w6907;
assign w6910 = A_357 & ~w6904;
assign w6911 = ~w6905 & w6910;
assign w6912 = ~A_357 & ~w6906;
assign w6913 = ~w6911 & ~w6912;
assign w6914 = A_360 & ~w6899;
assign w6915 = ~w6900 & w6914;
assign w6916 = ~A_360 & ~w6901;
assign w6917 = ~w6915 & ~w6916;
assign w6918 = ~w6913 & ~w6917;
assign w6919 = w6918 & w6920;
assign w6920 = ~w6908 & ~w6909;
assign w6921 = ~w6918 & ~w6920;
assign w6922 = ~w6919 & ~w6921;
assign w6923 = ~w6913 & w6917;
assign w6924 = w6913 & ~w6917;
assign w6925 = ~w6923 & ~w6924;
assign w6926 = w6918 & ~w6920;
assign w6927 = ~w6902 & ~w6907;
assign w6928 = ~w6926 & ~w6927;
assign w6929 = ~w6925 & ~w6928;
assign w6930 = ~w6922 & ~w6929;
assign w6931 = ~w6922 & ~w6928;
assign w6932 = A_364 & A_365;
assign w6933 = A_364 & ~A_365;
assign w6934 = ~A_364 & A_365;
assign w6935 = ~w6933 & ~w6934;
assign w6936 = (~w6932 & w6935) | (~w6932 & w12802) | (w6935 & w12802);
assign w6937 = A_361 & A_362;
assign w6938 = A_361 & ~A_362;
assign w6939 = ~A_361 & A_362;
assign w6940 = ~w6938 & ~w6939;
assign w6941 = (~w6937 & w6940) | (~w6937 & w12803) | (w6940 & w12803);
assign w6942 = ~w6936 & w6941;
assign w6943 = w6936 & ~w6941;
assign w6944 = ~w6942 & ~w6943;
assign w6945 = A_363 & ~w6938;
assign w6946 = ~w6939 & w6945;
assign w6947 = ~A_363 & ~w6940;
assign w6948 = ~w6946 & ~w6947;
assign w6949 = A_366 & ~w6933;
assign w6950 = ~w6934 & w6949;
assign w6951 = ~A_366 & ~w6935;
assign w6952 = ~w6950 & ~w6951;
assign w6953 = ~w6948 & ~w6952;
assign w6954 = ~w6944 & w6953;
assign w6955 = ~w6936 & ~w6941;
assign w6956 = ~w6954 & ~w6955;
assign w6957 = w6953 & w6944;
assign w6958 = ~w6944 & ~w6953;
assign w6959 = ~w6957 & ~w6958;
assign w6960 = ~w6956 & ~w6959;
assign w6961 = ~w6948 & w6952;
assign w6962 = w6948 & ~w6952;
assign w6963 = ~w6961 & ~w6962;
assign w6964 = ~w6925 & ~w6963;
assign w6965 = ~w6960 & w6964;
assign w6966 = ~w6931 & w6965;
assign w6967 = ~w6956 & ~w6963;
assign w6968 = ~w6959 & ~w6967;
assign w6969 = ~w6966 & ~w6968;
assign w6970 = ~w6959 & w6964;
assign w6971 = ~w6960 & w6970;
assign w6972 = ~w6931 & ~w6967;
assign w6973 = w6971 & w6972;
assign w6974 = (w6930 & w6969) | (w6930 & w13014) | (w6969 & w13014);
assign w6975 = ~w6966 & w6968;
assign w6976 = w6966 & ~w6968;
assign w6977 = ~w6975 & ~w6976;
assign w6978 = ~w6930 & ~w6977;
assign w6979 = ~w6960 & ~w6963;
assign w6980 = ~w6925 & ~w6931;
assign w6981 = ~w6979 & w6980;
assign w6982 = w6979 & ~w6980;
assign w6983 = ~w6981 & ~w6982;
assign w6984 = ~w6878 & ~w6881;
assign w6985 = ~w6843 & ~w6849;
assign w6986 = ~w6984 & w6985;
assign w6987 = w6984 & ~w6985;
assign w6988 = ~w6986 & ~w6987;
assign w6989 = ~w6983 & ~w6988;
assign w6990 = ~w6978 & w13015;
assign w6991 = (w6989 & w6978) | (w6989 & w13016) | (w6978 & w13016);
assign w6992 = ~w6990 & ~w6991;
assign w6993 = ~w6897 & ~w6992;
assign w6994 = ~w6978 & w13017;
assign w6995 = (~w6989 & w6978) | (~w6989 & w13400) | (w6978 & w13400);
assign w6996 = (w6897 & w6995) | (w6897 & w13018) | (w6995 & w13018);
assign w6997 = ~w6983 & w6988;
assign w6998 = w6983 & ~w6988;
assign w6999 = ~w6997 & ~w6998;
assign w7000 = ~w6718 & w6787;
assign w7001 = w6718 & ~w6787;
assign w7002 = ~w7000 & ~w7001;
assign w7003 = ~w6999 & ~w7002;
assign w7004 = ~w7003 & ~w6996;
assign w7005 = ~w6993 & w7004;
assign w7006 = ~w6993 & ~w6996;
assign w7007 = w7003 & ~w7006;
assign w7008 = (~w6815 & w7007) | (~w6815 & w13401) | (w7007 & w13401);
assign w7009 = w7003 & ~w6996;
assign w7010 = ~w6993 & w7009;
assign w7011 = ~w7003 & ~w7006;
assign w7012 = ~w7010 & ~w7011;
assign w7013 = (w6815 & w7011) | (w6815 & w13878) | (w7011 & w13878);
assign w7014 = ~w6999 & w7002;
assign w7015 = w6999 & ~w7002;
assign w7016 = ~w7014 & ~w7015;
assign w7017 = ~A_313 & A_314;
assign w7018 = A_313 & ~A_314;
assign w7019 = A_315 & ~w7018;
assign w7020 = ~w7017 & w7019;
assign w7021 = ~w7017 & ~w7018;
assign w7022 = ~A_315 & ~w7021;
assign w7023 = ~w7020 & ~w7022;
assign w7024 = ~A_316 & A_317;
assign w7025 = A_316 & ~A_317;
assign w7026 = A_318 & ~w7025;
assign w7027 = ~w7024 & w7026;
assign w7028 = ~w7024 & ~w7025;
assign w7029 = ~A_318 & ~w7028;
assign w7030 = ~w7027 & ~w7029;
assign w7031 = ~w7023 & w7030;
assign w7032 = w7023 & ~w7030;
assign w7033 = ~w7031 & ~w7032;
assign w7034 = A_316 & A_317;
assign w7035 = (~w7034 & w7028) | (~w7034 & w12804) | (w7028 & w12804);
assign w7036 = A_313 & A_314;
assign w7037 = (~w7036 & w7021) | (~w7036 & w12805) | (w7021 & w12805);
assign w7038 = ~w7035 & w7037;
assign w7039 = w7035 & ~w7037;
assign w7040 = ~w7038 & ~w7039;
assign w7041 = ~w7023 & ~w7030;
assign w7042 = ~w7040 & w7041;
assign w7043 = ~w7035 & ~w7037;
assign w7044 = ~w7042 & ~w7043;
assign w7045 = w7041 & w7040;
assign w7046 = ~w7040 & ~w7041;
assign w7047 = ~w7045 & ~w7046;
assign w7048 = ~w7044 & ~w7047;
assign w7049 = ~w7033 & ~w7048;
assign w7050 = ~A_307 & A_308;
assign w7051 = A_307 & ~A_308;
assign w7052 = A_309 & ~w7051;
assign w7053 = ~w7050 & w7052;
assign w7054 = ~w7050 & ~w7051;
assign w7055 = ~A_309 & ~w7054;
assign w7056 = ~w7053 & ~w7055;
assign w7057 = ~A_310 & A_311;
assign w7058 = A_310 & ~A_311;
assign w7059 = A_312 & ~w7058;
assign w7060 = ~w7057 & w7059;
assign w7061 = ~w7057 & ~w7058;
assign w7062 = ~A_312 & ~w7061;
assign w7063 = ~w7060 & ~w7062;
assign w7064 = ~w7056 & w7063;
assign w7065 = w7056 & ~w7063;
assign w7066 = ~w7064 & ~w7065;
assign w7067 = A_310 & A_311;
assign w7068 = (~w7067 & w7061) | (~w7067 & w12806) | (w7061 & w12806);
assign w7069 = A_307 & A_308;
assign w7070 = (~w7069 & w7054) | (~w7069 & w12807) | (w7054 & w12807);
assign w7071 = ~w7068 & w7070;
assign w7072 = w7068 & ~w7070;
assign w7073 = ~w7071 & ~w7072;
assign w7074 = ~w7056 & ~w7063;
assign w7075 = ~w7073 & w7074;
assign w7076 = ~w7068 & ~w7070;
assign w7077 = ~w7075 & ~w7076;
assign w7078 = w7074 & w7073;
assign w7079 = ~w7073 & ~w7074;
assign w7080 = ~w7078 & ~w7079;
assign w7081 = ~w7077 & ~w7080;
assign w7082 = ~w7066 & ~w7081;
assign w7083 = ~w7049 & w7082;
assign w7084 = w7049 & ~w7082;
assign w7085 = ~w7083 & ~w7084;
assign w7086 = ~A_301 & A_302;
assign w7087 = A_301 & ~A_302;
assign w7088 = A_303 & ~w7087;
assign w7089 = ~w7086 & w7088;
assign w7090 = ~w7086 & ~w7087;
assign w7091 = ~A_303 & ~w7090;
assign w7092 = ~w7089 & ~w7091;
assign w7093 = ~A_304 & A_305;
assign w7094 = A_304 & ~A_305;
assign w7095 = A_306 & ~w7094;
assign w7096 = ~w7093 & w7095;
assign w7097 = ~w7093 & ~w7094;
assign w7098 = ~A_306 & ~w7097;
assign w7099 = ~w7096 & ~w7098;
assign w7100 = ~w7092 & w7099;
assign w7101 = w7092 & ~w7099;
assign w7102 = ~w7100 & ~w7101;
assign w7103 = A_304 & A_305;
assign w7104 = (~w7103 & w7097) | (~w7103 & w12808) | (w7097 & w12808);
assign w7105 = A_301 & A_302;
assign w7106 = (~w7105 & w7090) | (~w7105 & w12809) | (w7090 & w12809);
assign w7107 = ~w7104 & w7106;
assign w7108 = w7104 & ~w7106;
assign w7109 = ~w7107 & ~w7108;
assign w7110 = ~w7092 & ~w7099;
assign w7111 = ~w7109 & w7110;
assign w7112 = ~w7104 & ~w7106;
assign w7113 = ~w7111 & ~w7112;
assign w7114 = w7110 & w7109;
assign w7115 = ~w7109 & ~w7110;
assign w7116 = ~w7114 & ~w7115;
assign w7117 = ~w7113 & ~w7116;
assign w7118 = ~w7102 & ~w7117;
assign w7119 = ~A_295 & A_296;
assign w7120 = A_295 & ~A_296;
assign w7121 = A_297 & ~w7120;
assign w7122 = ~w7119 & w7121;
assign w7123 = ~w7119 & ~w7120;
assign w7124 = ~A_297 & ~w7123;
assign w7125 = ~w7122 & ~w7124;
assign w7126 = ~A_298 & A_299;
assign w7127 = A_298 & ~A_299;
assign w7128 = A_300 & ~w7127;
assign w7129 = ~w7126 & w7128;
assign w7130 = ~w7126 & ~w7127;
assign w7131 = ~A_300 & ~w7130;
assign w7132 = ~w7129 & ~w7131;
assign w7133 = ~w7125 & w7132;
assign w7134 = w7125 & ~w7132;
assign w7135 = ~w7133 & ~w7134;
assign w7136 = A_298 & A_299;
assign w7137 = (~w7136 & w7130) | (~w7136 & w12810) | (w7130 & w12810);
assign w7138 = A_295 & A_296;
assign w7139 = (~w7138 & w7123) | (~w7138 & w12811) | (w7123 & w12811);
assign w7140 = ~w7137 & w7139;
assign w7141 = w7137 & ~w7139;
assign w7142 = ~w7140 & ~w7141;
assign w7143 = ~w7125 & ~w7132;
assign w7144 = ~w7142 & w7143;
assign w7145 = ~w7137 & ~w7139;
assign w7146 = ~w7144 & ~w7145;
assign w7147 = w7143 & w7142;
assign w7148 = ~w7142 & ~w7143;
assign w7149 = ~w7147 & ~w7148;
assign w7150 = ~w7146 & ~w7149;
assign w7151 = ~w7135 & ~w7150;
assign w7152 = ~w7118 & w7151;
assign w7153 = w7118 & ~w7151;
assign w7154 = ~w7152 & ~w7153;
assign w7155 = ~w7085 & w7154;
assign w7156 = w7085 & ~w7154;
assign w7157 = ~w7155 & ~w7156;
assign w7158 = ~A_289 & A_290;
assign w7159 = A_289 & ~A_290;
assign w7160 = A_291 & ~w7159;
assign w7161 = ~w7158 & w7160;
assign w7162 = ~w7158 & ~w7159;
assign w7163 = ~A_291 & ~w7162;
assign w7164 = ~w7161 & ~w7163;
assign w7165 = ~A_292 & A_293;
assign w7166 = A_292 & ~A_293;
assign w7167 = A_294 & ~w7166;
assign w7168 = ~w7165 & w7167;
assign w7169 = ~w7165 & ~w7166;
assign w7170 = ~A_294 & ~w7169;
assign w7171 = ~w7168 & ~w7170;
assign w7172 = ~w7164 & w7171;
assign w7173 = w7164 & ~w7171;
assign w7174 = ~w7172 & ~w7173;
assign w7175 = A_292 & A_293;
assign w7176 = (~w7175 & w7169) | (~w7175 & w12812) | (w7169 & w12812);
assign w7177 = A_289 & A_290;
assign w7178 = (~w7177 & w7162) | (~w7177 & w12813) | (w7162 & w12813);
assign w7179 = ~w7176 & w7178;
assign w7180 = w7176 & ~w7178;
assign w7181 = ~w7179 & ~w7180;
assign w7182 = ~w7164 & ~w7171;
assign w7183 = ~w7181 & w7182;
assign w7184 = ~w7176 & ~w7178;
assign w7185 = ~w7183 & ~w7184;
assign w7186 = w7182 & w7181;
assign w7187 = ~w7181 & ~w7182;
assign w7188 = ~w7186 & ~w7187;
assign w7189 = ~w7185 & ~w7188;
assign w7190 = ~w7174 & ~w7189;
assign w7191 = ~A_283 & A_284;
assign w7192 = A_283 & ~A_284;
assign w7193 = A_285 & ~w7192;
assign w7194 = ~w7191 & w7193;
assign w7195 = ~w7191 & ~w7192;
assign w7196 = ~A_285 & ~w7195;
assign w7197 = ~w7194 & ~w7196;
assign w7198 = ~A_286 & A_287;
assign w7199 = A_286 & ~A_287;
assign w7200 = A_288 & ~w7199;
assign w7201 = ~w7198 & w7200;
assign w7202 = ~w7198 & ~w7199;
assign w7203 = ~A_288 & ~w7202;
assign w7204 = ~w7201 & ~w7203;
assign w7205 = ~w7197 & w7204;
assign w7206 = w7197 & ~w7204;
assign w7207 = ~w7205 & ~w7206;
assign w7208 = A_286 & A_287;
assign w7209 = (~w7208 & w7202) | (~w7208 & w12814) | (w7202 & w12814);
assign w7210 = A_283 & A_284;
assign w7211 = (~w7210 & w7195) | (~w7210 & w12815) | (w7195 & w12815);
assign w7212 = ~w7209 & w7211;
assign w7213 = w7209 & ~w7211;
assign w7214 = ~w7212 & ~w7213;
assign w7215 = ~w7197 & ~w7204;
assign w7216 = ~w7214 & w7215;
assign w7217 = ~w7209 & ~w7211;
assign w7218 = ~w7216 & ~w7217;
assign w7219 = w7215 & w7214;
assign w7220 = ~w7214 & ~w7215;
assign w7221 = ~w7219 & ~w7220;
assign w7222 = ~w7218 & ~w7221;
assign w7223 = ~w7207 & ~w7222;
assign w7224 = ~w7190 & w7223;
assign w7225 = w7190 & ~w7223;
assign w7226 = ~w7224 & ~w7225;
assign w7227 = ~A_277 & A_278;
assign w7228 = A_277 & ~A_278;
assign w7229 = A_279 & ~w7228;
assign w7230 = ~w7227 & w7229;
assign w7231 = ~w7227 & ~w7228;
assign w7232 = ~A_279 & ~w7231;
assign w7233 = ~w7230 & ~w7232;
assign w7234 = ~A_280 & A_281;
assign w7235 = A_280 & ~A_281;
assign w7236 = A_282 & ~w7235;
assign w7237 = ~w7234 & w7236;
assign w7238 = ~w7234 & ~w7235;
assign w7239 = ~A_282 & ~w7238;
assign w7240 = ~w7237 & ~w7239;
assign w7241 = ~w7233 & w7240;
assign w7242 = w7233 & ~w7240;
assign w7243 = ~w7241 & ~w7242;
assign w7244 = A_280 & A_281;
assign w7245 = (~w7244 & w7238) | (~w7244 & w12816) | (w7238 & w12816);
assign w7246 = A_277 & A_278;
assign w7247 = (~w7246 & w7231) | (~w7246 & w12817) | (w7231 & w12817);
assign w7248 = ~w7245 & w7247;
assign w7249 = w7245 & ~w7247;
assign w7250 = ~w7248 & ~w7249;
assign w7251 = ~w7233 & ~w7240;
assign w7252 = ~w7250 & w7251;
assign w7253 = ~w7245 & ~w7247;
assign w7254 = ~w7252 & ~w7253;
assign w7255 = w7251 & w7250;
assign w7256 = ~w7250 & ~w7251;
assign w7257 = ~w7255 & ~w7256;
assign w7258 = ~w7254 & ~w7257;
assign w7259 = ~w7243 & ~w7258;
assign w7260 = ~A_271 & A_272;
assign w7261 = A_271 & ~A_272;
assign w7262 = A_273 & ~w7261;
assign w7263 = ~w7260 & w7262;
assign w7264 = ~w7260 & ~w7261;
assign w7265 = ~A_273 & ~w7264;
assign w7266 = ~w7263 & ~w7265;
assign w7267 = ~A_274 & A_275;
assign w7268 = A_274 & ~A_275;
assign w7269 = A_276 & ~w7268;
assign w7270 = ~w7267 & w7269;
assign w7271 = ~w7267 & ~w7268;
assign w7272 = ~A_276 & ~w7271;
assign w7273 = ~w7270 & ~w7272;
assign w7274 = ~w7266 & w7273;
assign w7275 = w7266 & ~w7273;
assign w7276 = ~w7274 & ~w7275;
assign w7277 = A_274 & A_275;
assign w7278 = (~w7277 & w7271) | (~w7277 & w12818) | (w7271 & w12818);
assign w7279 = A_271 & A_272;
assign w7280 = (~w7279 & w7264) | (~w7279 & w12819) | (w7264 & w12819);
assign w7281 = ~w7278 & w7280;
assign w7282 = w7278 & ~w7280;
assign w7283 = ~w7281 & ~w7282;
assign w7284 = ~w7266 & ~w7273;
assign w7285 = ~w7283 & w7284;
assign w7286 = ~w7278 & ~w7280;
assign w7287 = ~w7285 & ~w7286;
assign w7288 = w7284 & w7283;
assign w7289 = ~w7283 & ~w7284;
assign w7290 = ~w7288 & ~w7289;
assign w7291 = ~w7287 & ~w7290;
assign w7292 = ~w7276 & ~w7291;
assign w7293 = ~w7259 & w7292;
assign w7294 = w7259 & ~w7292;
assign w7295 = ~w7293 & ~w7294;
assign w7296 = ~w7226 & w7295;
assign w7297 = w7226 & ~w7295;
assign w7298 = ~w7296 & ~w7297;
assign w7299 = ~w7157 & w7298;
assign w7300 = w7157 & ~w7298;
assign w7301 = ~w7299 & ~w7300;
assign w7302 = ~w7016 & ~w7301;
assign w7303 = (w7302 & w7012) | (w7302 & w13402) | (w7012 & w13402);
assign w7304 = ~w7008 & w7303;
assign w7305 = (~w7302 & w7013) | (~w7302 & w13403) | (w7013 & w13403);
assign w7306 = ~w7304 & ~w7305;
assign w7307 = ~w7135 & ~w7146;
assign w7308 = ~w7149 & ~w7307;
assign w7309 = ~w7102 & ~w7135;
assign w7310 = ~w7117 & w7309;
assign w7311 = ~w7150 & w7310;
assign w7312 = ~w7102 & ~w7113;
assign w7313 = ~w7116 & ~w7312;
assign w7314 = ~w7311 & w7313;
assign w7315 = w7311 & ~w7313;
assign w7316 = ~w7314 & ~w7315;
assign w7317 = ~w7308 & ~w7316;
assign w7318 = ~w7311 & ~w7313;
assign w7319 = ~w7116 & w7309;
assign w7320 = ~w7117 & w7319;
assign w7321 = ~w7150 & ~w7312;
assign w7322 = w7320 & w7321;
assign w7323 = (w7308 & w7318) | (w7308 & w13404) | (w7318 & w13404);
assign w7324 = ~w7317 & ~w7323;
assign w7325 = ~w7066 & ~w7077;
assign w7326 = ~w7080 & ~w7325;
assign w7327 = ~w7033 & ~w7066;
assign w7328 = ~w7048 & w7327;
assign w7329 = ~w7081 & w7328;
assign w7330 = ~w7033 & ~w7044;
assign w7331 = ~w7047 & ~w7330;
assign w7332 = ~w7329 & ~w7331;
assign w7333 = ~w7047 & w7327;
assign w7334 = ~w7048 & w7333;
assign w7335 = ~w7081 & ~w7330;
assign w7336 = w7334 & w7335;
assign w7337 = (w7326 & w7332) | (w7326 & w13019) | (w7332 & w13019);
assign w7338 = ~w7329 & w7331;
assign w7339 = w7329 & ~w7331;
assign w7340 = ~w7338 & ~w7339;
assign w7341 = ~w7326 & ~w7340;
assign w7342 = ~w7085 & ~w7154;
assign w7343 = ~w7341 & w13020;
assign w7344 = (w7342 & w7341) | (w7342 & w13021) | (w7341 & w13021);
assign w7345 = ~w7343 & ~w7344;
assign w7346 = ~w7324 & ~w7345;
assign w7347 = ~w7341 & w13022;
assign w7348 = (~w7342 & w7341) | (~w7342 & w13405) | (w7341 & w13405);
assign w7349 = (w7324 & w7348) | (w7324 & w13023) | (w7348 & w13023);
assign w7350 = ~w7157 & ~w7298;
assign w7351 = w7350 & ~w7349;
assign w7352 = ~w7346 & w7351;
assign w7353 = ~w7346 & ~w7349;
assign w7354 = ~w7350 & ~w7353;
assign w7355 = ~w7207 & ~w7218;
assign w7356 = ~w7221 & ~w7355;
assign w7357 = ~w7174 & ~w7207;
assign w7358 = ~w7189 & w7357;
assign w7359 = ~w7222 & w7358;
assign w7360 = ~w7174 & ~w7185;
assign w7361 = ~w7188 & ~w7360;
assign w7362 = ~w7359 & ~w7361;
assign w7363 = ~w7188 & w7357;
assign w7364 = ~w7189 & w7363;
assign w7365 = ~w7222 & ~w7360;
assign w7366 = w7364 & w7365;
assign w7367 = (w7356 & w7362) | (w7356 & w13024) | (w7362 & w13024);
assign w7368 = ~w7359 & w7361;
assign w7369 = w7359 & ~w7361;
assign w7370 = ~w7368 & ~w7369;
assign w7371 = ~w7356 & ~w7370;
assign w7372 = ~w7226 & ~w7295;
assign w7373 = ~w7371 & w13406;
assign w7374 = (~w7372 & w7371) | (~w7372 & w13407) | (w7371 & w13407);
assign w7375 = ~w7373 & ~w7374;
assign w7376 = ~w7276 & ~w7287;
assign w7377 = ~w7290 & ~w7376;
assign w7378 = ~w7243 & ~w7276;
assign w7379 = ~w7258 & w7378;
assign w7380 = ~w7291 & w7379;
assign w7381 = ~w7243 & ~w7254;
assign w7382 = ~w7257 & ~w7381;
assign w7383 = ~w7380 & w7382;
assign w7384 = w7380 & ~w7382;
assign w7385 = ~w7383 & ~w7384;
assign w7386 = ~w7377 & ~w7385;
assign w7387 = ~w7380 & ~w7382;
assign w7388 = ~w7257 & w7378;
assign w7389 = ~w7258 & w7388;
assign w7390 = ~w7291 & ~w7381;
assign w7391 = w7389 & w7390;
assign w7392 = (w7377 & w7387) | (w7377 & w13408) | (w7387 & w13408);
assign w7393 = ~w7386 & ~w7392;
assign w7394 = ~w7375 & w7393;
assign w7395 = ~w7371 & w13025;
assign w7396 = (w7372 & w7371) | (w7372 & w13409) | (w7371 & w13409);
assign w7397 = ~w7395 & ~w7396;
assign w7398 = ~w7393 & ~w7397;
assign w7399 = ~w7394 & ~w7398;
assign w7400 = (w7399 & w7354) | (w7399 & w13879) | (w7354 & w13879);
assign w7401 = ~w7350 & ~w7349;
assign w7402 = ~w7346 & w7401;
assign w7403 = w7350 & ~w7353;
assign w7404 = (~w7399 & w7403) | (~w7399 & w13880) | (w7403 & w13880);
assign w7405 = ~w7400 & ~w7404;
assign w7406 = ~w7306 & w7405;
assign w7407 = (~w7302 & w7012) | (~w7302 & w13410) | (w7012 & w13410);
assign w7408 = ~w7008 & w7407;
assign w7409 = (w7302 & w7013) | (w7302 & w13411) | (w7013 & w13411);
assign w7410 = ~w7408 & ~w7409;
assign w7411 = ~w7405 & ~w7410;
assign w7412 = ~w7406 & ~w7411;
assign w7413 = A_394 & A_395;
assign w7414 = A_394 & ~A_395;
assign w7415 = ~A_394 & A_395;
assign w7416 = ~w7414 & ~w7415;
assign w7417 = (~w7413 & w7416) | (~w7413 & w12820) | (w7416 & w12820);
assign w7418 = A_391 & A_392;
assign w7419 = A_391 & ~A_392;
assign w7420 = ~A_391 & A_392;
assign w7421 = ~w7419 & ~w7420;
assign w7422 = (~w7418 & w7421) | (~w7418 & w12821) | (w7421 & w12821);
assign w7423 = w7417 & ~w7422;
assign w7424 = ~w7417 & w7422;
assign w7425 = A_393 & ~w7419;
assign w7426 = ~w7420 & w7425;
assign w7427 = ~A_393 & ~w7421;
assign w7428 = ~w7426 & ~w7427;
assign w7429 = A_396 & ~w7414;
assign w7430 = ~w7415 & w7429;
assign w7431 = ~A_396 & ~w7416;
assign w7432 = ~w7430 & ~w7431;
assign w7433 = ~w7428 & ~w7432;
assign w7434 = w7433 & w7435;
assign w7435 = ~w7423 & ~w7424;
assign w7436 = ~w7433 & ~w7435;
assign w7437 = ~w7434 & ~w7436;
assign w7438 = ~w7428 & w7432;
assign w7439 = w7428 & ~w7432;
assign w7440 = ~w7438 & ~w7439;
assign w7441 = w7433 & ~w7435;
assign w7442 = ~w7417 & ~w7422;
assign w7443 = ~w7441 & ~w7442;
assign w7444 = ~w7440 & ~w7443;
assign w7445 = ~w7437 & ~w7444;
assign w7446 = ~w7437 & ~w7443;
assign w7447 = A_400 & A_401;
assign w7448 = A_400 & ~A_401;
assign w7449 = ~A_400 & A_401;
assign w7450 = ~w7448 & ~w7449;
assign w7451 = (~w7447 & w7450) | (~w7447 & w12822) | (w7450 & w12822);
assign w7452 = A_397 & A_398;
assign w7453 = A_397 & ~A_398;
assign w7454 = ~A_397 & A_398;
assign w7455 = ~w7453 & ~w7454;
assign w7456 = (~w7452 & w7455) | (~w7452 & w12823) | (w7455 & w12823);
assign w7457 = ~w7451 & w7456;
assign w7458 = w7451 & ~w7456;
assign w7459 = ~w7457 & ~w7458;
assign w7460 = A_399 & ~w7453;
assign w7461 = ~w7454 & w7460;
assign w7462 = ~A_399 & ~w7455;
assign w7463 = ~w7461 & ~w7462;
assign w7464 = A_402 & ~w7448;
assign w7465 = ~w7449 & w7464;
assign w7466 = ~A_402 & ~w7450;
assign w7467 = ~w7465 & ~w7466;
assign w7468 = ~w7463 & ~w7467;
assign w7469 = ~w7459 & w7468;
assign w7470 = ~w7451 & ~w7456;
assign w7471 = ~w7469 & ~w7470;
assign w7472 = w7468 & w7459;
assign w7473 = ~w7459 & ~w7468;
assign w7474 = ~w7472 & ~w7473;
assign w7475 = ~w7471 & ~w7474;
assign w7476 = ~w7463 & w7467;
assign w7477 = w7463 & ~w7467;
assign w7478 = ~w7476 & ~w7477;
assign w7479 = ~w7440 & ~w7478;
assign w7480 = ~w7475 & w7479;
assign w7481 = ~w7446 & w7480;
assign w7482 = ~w7471 & ~w7478;
assign w7483 = ~w7474 & ~w7482;
assign w7484 = ~w7481 & w7483;
assign w7485 = w7481 & ~w7483;
assign w7486 = ~w7484 & ~w7485;
assign w7487 = ~w7445 & ~w7486;
assign w7488 = ~w7481 & ~w7483;
assign w7489 = ~w7474 & w7479;
assign w7490 = ~w7475 & w7489;
assign w7491 = ~w7446 & ~w7482;
assign w7492 = w7490 & w7491;
assign w7493 = (w7445 & w7488) | (w7445 & w13412) | (w7488 & w13412);
assign w7494 = ~w7487 & ~w7493;
assign w7495 = A_406 & A_407;
assign w7496 = A_406 & ~A_407;
assign w7497 = ~A_406 & A_407;
assign w7498 = ~w7496 & ~w7497;
assign w7499 = (~w7495 & w7498) | (~w7495 & w12824) | (w7498 & w12824);
assign w7500 = A_403 & A_404;
assign w7501 = A_403 & ~A_404;
assign w7502 = ~A_403 & A_404;
assign w7503 = ~w7501 & ~w7502;
assign w7504 = (~w7500 & w7503) | (~w7500 & w12825) | (w7503 & w12825);
assign w7505 = w7499 & ~w7504;
assign w7506 = ~w7499 & w7504;
assign w7507 = A_405 & ~w7501;
assign w7508 = ~w7502 & w7507;
assign w7509 = ~A_405 & ~w7503;
assign w7510 = ~w7508 & ~w7509;
assign w7511 = A_408 & ~w7496;
assign w7512 = ~w7497 & w7511;
assign w7513 = ~A_408 & ~w7498;
assign w7514 = ~w7512 & ~w7513;
assign w7515 = ~w7510 & ~w7514;
assign w7516 = w7515 & w7517;
assign w7517 = ~w7505 & ~w7506;
assign w7518 = ~w7515 & ~w7517;
assign w7519 = ~w7516 & ~w7518;
assign w7520 = ~w7510 & w7514;
assign w7521 = w7510 & ~w7514;
assign w7522 = ~w7520 & ~w7521;
assign w7523 = w7515 & ~w7517;
assign w7524 = ~w7499 & ~w7504;
assign w7525 = ~w7523 & ~w7524;
assign w7526 = ~w7522 & ~w7525;
assign w7527 = ~w7519 & ~w7526;
assign w7528 = ~w7519 & ~w7525;
assign w7529 = A_412 & A_413;
assign w7530 = A_412 & ~A_413;
assign w7531 = ~A_412 & A_413;
assign w7532 = ~w7530 & ~w7531;
assign w7533 = (~w7529 & w7532) | (~w7529 & w12826) | (w7532 & w12826);
assign w7534 = A_409 & A_410;
assign w7535 = A_409 & ~A_410;
assign w7536 = ~A_409 & A_410;
assign w7537 = ~w7535 & ~w7536;
assign w7538 = (~w7534 & w7537) | (~w7534 & w12827) | (w7537 & w12827);
assign w7539 = ~w7533 & w7538;
assign w7540 = w7533 & ~w7538;
assign w7541 = ~w7539 & ~w7540;
assign w7542 = A_411 & ~w7535;
assign w7543 = ~w7536 & w7542;
assign w7544 = ~A_411 & ~w7537;
assign w7545 = ~w7543 & ~w7544;
assign w7546 = A_414 & ~w7530;
assign w7547 = ~w7531 & w7546;
assign w7548 = ~A_414 & ~w7532;
assign w7549 = ~w7547 & ~w7548;
assign w7550 = ~w7545 & ~w7549;
assign w7551 = ~w7541 & w7550;
assign w7552 = ~w7533 & ~w7538;
assign w7553 = ~w7551 & ~w7552;
assign w7554 = w7550 & w7541;
assign w7555 = ~w7541 & ~w7550;
assign w7556 = ~w7554 & ~w7555;
assign w7557 = ~w7553 & ~w7556;
assign w7558 = ~w7545 & w7549;
assign w7559 = w7545 & ~w7549;
assign w7560 = ~w7558 & ~w7559;
assign w7561 = ~w7522 & ~w7560;
assign w7562 = ~w7557 & w7561;
assign w7563 = ~w7528 & w7562;
assign w7564 = ~w7553 & ~w7560;
assign w7565 = ~w7556 & ~w7564;
assign w7566 = ~w7563 & ~w7565;
assign w7567 = ~w7556 & w7561;
assign w7568 = ~w7557 & w7567;
assign w7569 = ~w7528 & ~w7564;
assign w7570 = w7568 & w7569;
assign w7571 = (w7527 & w7566) | (w7527 & w13026) | (w7566 & w13026);
assign w7572 = ~w7563 & w7565;
assign w7573 = w7563 & ~w7565;
assign w7574 = ~w7572 & ~w7573;
assign w7575 = ~w7527 & ~w7574;
assign w7576 = ~w7557 & ~w7560;
assign w7577 = ~w7522 & ~w7528;
assign w7578 = ~w7576 & w7577;
assign w7579 = w7576 & ~w7577;
assign w7580 = ~w7578 & ~w7579;
assign w7581 = ~w7475 & ~w7478;
assign w7582 = ~w7440 & ~w7446;
assign w7583 = ~w7581 & w7582;
assign w7584 = w7581 & ~w7582;
assign w7585 = ~w7583 & ~w7584;
assign w7586 = ~w7580 & ~w7585;
assign w7587 = ~w7575 & w13027;
assign w7588 = (w7586 & w7575) | (w7586 & w13028) | (w7575 & w13028);
assign w7589 = ~w7587 & ~w7588;
assign w7590 = ~w7494 & ~w7589;
assign w7591 = ~w7575 & w13029;
assign w7592 = (~w7586 & w7575) | (~w7586 & w13413) | (w7575 & w13413);
assign w7593 = (w7494 & w7592) | (w7494 & w13030) | (w7592 & w13030);
assign w7594 = ~w7580 & w7585;
assign w7595 = w7580 & ~w7585;
assign w7596 = ~w7594 & ~w7595;
assign w7597 = ~A_385 & A_386;
assign w7598 = A_385 & ~A_386;
assign w7599 = A_387 & ~w7598;
assign w7600 = ~w7597 & w7599;
assign w7601 = ~w7597 & ~w7598;
assign w7602 = ~A_387 & ~w7601;
assign w7603 = ~w7600 & ~w7602;
assign w7604 = ~A_388 & A_389;
assign w7605 = A_388 & ~A_389;
assign w7606 = A_390 & ~w7605;
assign w7607 = ~w7604 & w7606;
assign w7608 = ~w7604 & ~w7605;
assign w7609 = ~A_390 & ~w7608;
assign w7610 = ~w7607 & ~w7609;
assign w7611 = ~w7603 & w7610;
assign w7612 = w7603 & ~w7610;
assign w7613 = ~w7611 & ~w7612;
assign w7614 = A_388 & A_389;
assign w7615 = (~w7614 & w7608) | (~w7614 & w12828) | (w7608 & w12828);
assign w7616 = A_385 & A_386;
assign w7617 = (~w7616 & w7601) | (~w7616 & w12829) | (w7601 & w12829);
assign w7618 = ~w7615 & w7617;
assign w7619 = w7615 & ~w7617;
assign w7620 = ~w7618 & ~w7619;
assign w7621 = ~w7603 & ~w7610;
assign w7622 = ~w7620 & w7621;
assign w7623 = ~w7615 & ~w7617;
assign w7624 = ~w7622 & ~w7623;
assign w7625 = w7621 & w7620;
assign w7626 = ~w7620 & ~w7621;
assign w7627 = ~w7625 & ~w7626;
assign w7628 = ~w7624 & ~w7627;
assign w7629 = ~w7613 & ~w7628;
assign w7630 = ~A_379 & A_380;
assign w7631 = A_379 & ~A_380;
assign w7632 = A_381 & ~w7631;
assign w7633 = ~w7630 & w7632;
assign w7634 = ~w7630 & ~w7631;
assign w7635 = ~A_381 & ~w7634;
assign w7636 = ~w7633 & ~w7635;
assign w7637 = ~A_382 & A_383;
assign w7638 = A_382 & ~A_383;
assign w7639 = A_384 & ~w7638;
assign w7640 = ~w7637 & w7639;
assign w7641 = ~w7637 & ~w7638;
assign w7642 = ~A_384 & ~w7641;
assign w7643 = ~w7640 & ~w7642;
assign w7644 = ~w7636 & w7643;
assign w7645 = w7636 & ~w7643;
assign w7646 = ~w7644 & ~w7645;
assign w7647 = A_382 & A_383;
assign w7648 = (~w7647 & w7641) | (~w7647 & w12830) | (w7641 & w12830);
assign w7649 = A_379 & A_380;
assign w7650 = (~w7649 & w7634) | (~w7649 & w12831) | (w7634 & w12831);
assign w7651 = ~w7648 & w7650;
assign w7652 = w7648 & ~w7650;
assign w7653 = ~w7651 & ~w7652;
assign w7654 = ~w7636 & ~w7643;
assign w7655 = ~w7653 & w7654;
assign w7656 = ~w7648 & ~w7650;
assign w7657 = ~w7655 & ~w7656;
assign w7658 = w7654 & w7653;
assign w7659 = ~w7653 & ~w7654;
assign w7660 = ~w7658 & ~w7659;
assign w7661 = ~w7657 & ~w7660;
assign w7662 = ~w7646 & ~w7661;
assign w7663 = ~w7629 & w7662;
assign w7664 = w7629 & ~w7662;
assign w7665 = ~w7663 & ~w7664;
assign w7666 = ~A_373 & A_374;
assign w7667 = A_373 & ~A_374;
assign w7668 = A_375 & ~w7667;
assign w7669 = ~w7666 & w7668;
assign w7670 = ~w7666 & ~w7667;
assign w7671 = ~A_375 & ~w7670;
assign w7672 = ~w7669 & ~w7671;
assign w7673 = ~A_376 & A_377;
assign w7674 = A_376 & ~A_377;
assign w7675 = A_378 & ~w7674;
assign w7676 = ~w7673 & w7675;
assign w7677 = ~w7673 & ~w7674;
assign w7678 = ~A_378 & ~w7677;
assign w7679 = ~w7676 & ~w7678;
assign w7680 = ~w7672 & w7679;
assign w7681 = w7672 & ~w7679;
assign w7682 = ~w7680 & ~w7681;
assign w7683 = A_376 & A_377;
assign w7684 = (~w7683 & w7677) | (~w7683 & w12832) | (w7677 & w12832);
assign w7685 = A_373 & A_374;
assign w7686 = (~w7685 & w7670) | (~w7685 & w12833) | (w7670 & w12833);
assign w7687 = ~w7684 & w7686;
assign w7688 = w7684 & ~w7686;
assign w7689 = ~w7687 & ~w7688;
assign w7690 = ~w7672 & ~w7679;
assign w7691 = ~w7689 & w7690;
assign w7692 = ~w7684 & ~w7686;
assign w7693 = ~w7691 & ~w7692;
assign w7694 = w7690 & w7689;
assign w7695 = ~w7689 & ~w7690;
assign w7696 = ~w7694 & ~w7695;
assign w7697 = ~w7693 & ~w7696;
assign w7698 = ~w7682 & ~w7697;
assign w7699 = ~A_367 & A_368;
assign w7700 = A_367 & ~A_368;
assign w7701 = A_369 & ~w7700;
assign w7702 = ~w7699 & w7701;
assign w7703 = ~w7699 & ~w7700;
assign w7704 = ~A_369 & ~w7703;
assign w7705 = ~w7702 & ~w7704;
assign w7706 = ~A_370 & A_371;
assign w7707 = A_370 & ~A_371;
assign w7708 = A_372 & ~w7707;
assign w7709 = ~w7706 & w7708;
assign w7710 = ~w7706 & ~w7707;
assign w7711 = ~A_372 & ~w7710;
assign w7712 = ~w7709 & ~w7711;
assign w7713 = ~w7705 & w7712;
assign w7714 = w7705 & ~w7712;
assign w7715 = ~w7713 & ~w7714;
assign w7716 = A_370 & A_371;
assign w7717 = (~w7716 & w7710) | (~w7716 & w12834) | (w7710 & w12834);
assign w7718 = A_367 & A_368;
assign w7719 = (~w7718 & w7703) | (~w7718 & w12835) | (w7703 & w12835);
assign w7720 = ~w7717 & w7719;
assign w7721 = w7717 & ~w7719;
assign w7722 = ~w7720 & ~w7721;
assign w7723 = ~w7705 & ~w7712;
assign w7724 = ~w7722 & w7723;
assign w7725 = ~w7717 & ~w7719;
assign w7726 = ~w7724 & ~w7725;
assign w7727 = w7723 & w7722;
assign w7728 = ~w7722 & ~w7723;
assign w7729 = ~w7727 & ~w7728;
assign w7730 = ~w7726 & ~w7729;
assign w7731 = ~w7715 & ~w7730;
assign w7732 = ~w7698 & w7731;
assign w7733 = w7698 & ~w7731;
assign w7734 = ~w7732 & ~w7733;
assign w7735 = ~w7665 & w7734;
assign w7736 = w7665 & ~w7734;
assign w7737 = ~w7735 & ~w7736;
assign w7738 = ~w7596 & ~w7737;
assign w7739 = w7738 & ~w7593;
assign w7740 = ~w7590 & w7739;
assign w7741 = ~w7590 & ~w7593;
assign w7742 = ~w7738 & ~w7741;
assign w7743 = ~w7646 & ~w7657;
assign w7744 = ~w7660 & ~w7743;
assign w7745 = ~w7613 & ~w7646;
assign w7746 = ~w7628 & w7745;
assign w7747 = ~w7661 & w7746;
assign w7748 = ~w7613 & ~w7624;
assign w7749 = ~w7627 & ~w7748;
assign w7750 = ~w7747 & ~w7749;
assign w7751 = ~w7627 & w7745;
assign w7752 = ~w7628 & w7751;
assign w7753 = ~w7661 & ~w7748;
assign w7754 = w7752 & w7753;
assign w7755 = (w7744 & w7750) | (w7744 & w13031) | (w7750 & w13031);
assign w7756 = ~w7747 & w7749;
assign w7757 = w7747 & ~w7749;
assign w7758 = ~w7756 & ~w7757;
assign w7759 = ~w7744 & ~w7758;
assign w7760 = ~w7665 & ~w7734;
assign w7761 = ~w7759 & w13414;
assign w7762 = (~w7760 & w7759) | (~w7760 & w13415) | (w7759 & w13415);
assign w7763 = ~w7761 & ~w7762;
assign w7764 = ~w7715 & ~w7726;
assign w7765 = ~w7729 & ~w7764;
assign w7766 = ~w7682 & ~w7715;
assign w7767 = ~w7697 & w7766;
assign w7768 = ~w7730 & w7767;
assign w7769 = ~w7682 & ~w7693;
assign w7770 = ~w7696 & ~w7769;
assign w7771 = ~w7768 & w7770;
assign w7772 = w7768 & ~w7770;
assign w7773 = ~w7771 & ~w7772;
assign w7774 = ~w7765 & ~w7773;
assign w7775 = ~w7768 & ~w7770;
assign w7776 = ~w7696 & w7766;
assign w7777 = ~w7697 & w7776;
assign w7778 = ~w7730 & ~w7769;
assign w7779 = w7777 & w7778;
assign w7780 = (w7765 & w7775) | (w7765 & w13416) | (w7775 & w13416);
assign w7781 = ~w7774 & ~w7780;
assign w7782 = ~w7763 & w7781;
assign w7783 = ~w7759 & w13032;
assign w7784 = (w7760 & w7759) | (w7760 & w13417) | (w7759 & w13417);
assign w7785 = ~w7783 & ~w7784;
assign w7786 = ~w7781 & ~w7785;
assign w7787 = ~w7782 & ~w7786;
assign w7788 = (w7787 & w7742) | (w7787 & w13418) | (w7742 & w13418);
assign w7789 = ~w7738 & ~w7593;
assign w7790 = ~w7590 & w7789;
assign w7791 = w7738 & ~w7741;
assign w7792 = (~w7787 & w7791) | (~w7787 & w13538) | (w7791 & w13538);
assign w7793 = ~w7788 & ~w7792;
assign w7794 = A_430 & A_431;
assign w7795 = A_430 & ~A_431;
assign w7796 = ~A_430 & A_431;
assign w7797 = ~w7795 & ~w7796;
assign w7798 = (~w7794 & w7797) | (~w7794 & w12836) | (w7797 & w12836);
assign w7799 = A_427 & A_428;
assign w7800 = A_427 & ~A_428;
assign w7801 = ~A_427 & A_428;
assign w7802 = ~w7800 & ~w7801;
assign w7803 = (~w7799 & w7802) | (~w7799 & w12837) | (w7802 & w12837);
assign w7804 = w7798 & ~w7803;
assign w7805 = ~w7798 & w7803;
assign w7806 = A_429 & ~w7800;
assign w7807 = ~w7801 & w7806;
assign w7808 = ~A_429 & ~w7802;
assign w7809 = ~w7807 & ~w7808;
assign w7810 = A_432 & ~w7795;
assign w7811 = ~w7796 & w7810;
assign w7812 = ~A_432 & ~w7797;
assign w7813 = ~w7811 & ~w7812;
assign w7814 = ~w7809 & ~w7813;
assign w7815 = w7814 & w7816;
assign w7816 = ~w7804 & ~w7805;
assign w7817 = ~w7814 & ~w7816;
assign w7818 = ~w7815 & ~w7817;
assign w7819 = ~w7809 & w7813;
assign w7820 = w7809 & ~w7813;
assign w7821 = ~w7819 & ~w7820;
assign w7822 = w7814 & ~w7816;
assign w7823 = ~w7798 & ~w7803;
assign w7824 = ~w7822 & ~w7823;
assign w7825 = ~w7821 & ~w7824;
assign w7826 = ~w7818 & ~w7825;
assign w7827 = ~w7818 & ~w7824;
assign w7828 = A_436 & A_437;
assign w7829 = A_436 & ~A_437;
assign w7830 = ~A_436 & A_437;
assign w7831 = ~w7829 & ~w7830;
assign w7832 = (~w7828 & w7831) | (~w7828 & w12838) | (w7831 & w12838);
assign w7833 = A_433 & A_434;
assign w7834 = A_433 & ~A_434;
assign w7835 = ~A_433 & A_434;
assign w7836 = ~w7834 & ~w7835;
assign w7837 = (~w7833 & w7836) | (~w7833 & w12839) | (w7836 & w12839);
assign w7838 = ~w7832 & w7837;
assign w7839 = w7832 & ~w7837;
assign w7840 = ~w7838 & ~w7839;
assign w7841 = A_435 & ~w7834;
assign w7842 = ~w7835 & w7841;
assign w7843 = ~A_435 & ~w7836;
assign w7844 = ~w7842 & ~w7843;
assign w7845 = A_438 & ~w7829;
assign w7846 = ~w7830 & w7845;
assign w7847 = ~A_438 & ~w7831;
assign w7848 = ~w7846 & ~w7847;
assign w7849 = ~w7844 & ~w7848;
assign w7850 = ~w7840 & w7849;
assign w7851 = ~w7832 & ~w7837;
assign w7852 = ~w7850 & ~w7851;
assign w7853 = w7849 & w7840;
assign w7854 = ~w7840 & ~w7849;
assign w7855 = ~w7853 & ~w7854;
assign w7856 = ~w7852 & ~w7855;
assign w7857 = ~w7844 & w7848;
assign w7858 = w7844 & ~w7848;
assign w7859 = ~w7857 & ~w7858;
assign w7860 = ~w7821 & ~w7859;
assign w7861 = ~w7856 & w7860;
assign w7862 = ~w7827 & w7861;
assign w7863 = ~w7852 & ~w7859;
assign w7864 = ~w7855 & ~w7863;
assign w7865 = ~w7862 & ~w7864;
assign w7866 = ~w7855 & w7860;
assign w7867 = ~w7856 & w7866;
assign w7868 = ~w7827 & ~w7863;
assign w7869 = w7867 & w7868;
assign w7870 = (w7826 & w7865) | (w7826 & w13033) | (w7865 & w13033);
assign w7871 = ~w7862 & w7864;
assign w7872 = w7862 & ~w7864;
assign w7873 = ~w7871 & ~w7872;
assign w7874 = ~w7826 & ~w7873;
assign w7875 = ~w7856 & ~w7859;
assign w7876 = ~w7821 & ~w7827;
assign w7877 = ~w7875 & w7876;
assign w7878 = w7875 & ~w7876;
assign w7879 = ~w7877 & ~w7878;
assign w7880 = ~A_421 & A_422;
assign w7881 = A_421 & ~A_422;
assign w7882 = A_423 & ~w7881;
assign w7883 = ~w7880 & w7882;
assign w7884 = ~w7880 & ~w7881;
assign w7885 = ~A_423 & ~w7884;
assign w7886 = ~w7883 & ~w7885;
assign w7887 = ~A_424 & A_425;
assign w7888 = A_424 & ~A_425;
assign w7889 = A_426 & ~w7888;
assign w7890 = ~w7887 & w7889;
assign w7891 = ~w7887 & ~w7888;
assign w7892 = ~A_426 & ~w7891;
assign w7893 = ~w7890 & ~w7892;
assign w7894 = ~w7886 & w7893;
assign w7895 = w7886 & ~w7893;
assign w7896 = ~w7894 & ~w7895;
assign w7897 = A_424 & A_425;
assign w7898 = (~w7897 & w7891) | (~w7897 & w12840) | (w7891 & w12840);
assign w7899 = A_421 & A_422;
assign w7900 = (~w7899 & w7884) | (~w7899 & w12841) | (w7884 & w12841);
assign w7901 = ~w7898 & w7900;
assign w7902 = w7898 & ~w7900;
assign w7903 = ~w7901 & ~w7902;
assign w7904 = ~w7886 & ~w7893;
assign w7905 = ~w7903 & w7904;
assign w7906 = ~w7898 & ~w7900;
assign w7907 = ~w7905 & ~w7906;
assign w7908 = w7904 & w7903;
assign w7909 = ~w7903 & ~w7904;
assign w7910 = ~w7908 & ~w7909;
assign w7911 = ~w7907 & ~w7910;
assign w7912 = ~w7896 & ~w7911;
assign w7913 = ~A_415 & A_416;
assign w7914 = A_415 & ~A_416;
assign w7915 = A_417 & ~w7914;
assign w7916 = ~w7913 & w7915;
assign w7917 = ~w7913 & ~w7914;
assign w7918 = ~A_417 & ~w7917;
assign w7919 = ~w7916 & ~w7918;
assign w7920 = ~A_418 & A_419;
assign w7921 = A_418 & ~A_419;
assign w7922 = A_420 & ~w7921;
assign w7923 = ~w7920 & w7922;
assign w7924 = ~w7920 & ~w7921;
assign w7925 = ~A_420 & ~w7924;
assign w7926 = ~w7923 & ~w7925;
assign w7927 = ~w7919 & w7926;
assign w7928 = w7919 & ~w7926;
assign w7929 = ~w7927 & ~w7928;
assign w7930 = A_418 & A_419;
assign w7931 = (~w7930 & w7924) | (~w7930 & w12842) | (w7924 & w12842);
assign w7932 = A_415 & A_416;
assign w7933 = (~w7932 & w7917) | (~w7932 & w12843) | (w7917 & w12843);
assign w7934 = ~w7931 & w7933;
assign w7935 = w7931 & ~w7933;
assign w7936 = ~w7934 & ~w7935;
assign w7937 = ~w7919 & ~w7926;
assign w7938 = ~w7936 & w7937;
assign w7939 = ~w7931 & ~w7933;
assign w7940 = ~w7938 & ~w7939;
assign w7941 = w7937 & w7936;
assign w7942 = ~w7936 & ~w7937;
assign w7943 = ~w7941 & ~w7942;
assign w7944 = ~w7940 & ~w7943;
assign w7945 = ~w7929 & ~w7944;
assign w7946 = ~w7912 & w7945;
assign w7947 = w7912 & ~w7945;
assign w7948 = ~w7946 & ~w7947;
assign w7949 = ~w7879 & ~w7948;
assign w7950 = ~w7874 & w13034;
assign w7951 = (~w7949 & w7874) | (~w7949 & w13035) | (w7874 & w13035);
assign w7952 = ~w7950 & ~w7951;
assign w7953 = ~w7929 & ~w7940;
assign w7954 = ~w7943 & ~w7953;
assign w7955 = ~w7896 & ~w7929;
assign w7956 = ~w7911 & w7955;
assign w7957 = ~w7944 & w7956;
assign w7958 = ~w7896 & ~w7907;
assign w7959 = ~w7910 & ~w7958;
assign w7960 = ~w7957 & w7959;
assign w7961 = w7957 & ~w7959;
assign w7962 = ~w7960 & ~w7961;
assign w7963 = ~w7954 & ~w7962;
assign w7964 = ~w7957 & ~w7959;
assign w7965 = ~w7910 & w7955;
assign w7966 = ~w7911 & w7965;
assign w7967 = ~w7944 & ~w7958;
assign w7968 = w7966 & w7967;
assign w7969 = (w7954 & w7964) | (w7954 & w13419) | (w7964 & w13419);
assign w7970 = ~w7963 & ~w7969;
assign w7971 = ~w7952 & w7970;
assign w7972 = ~w7874 & w13036;
assign w7973 = (w7949 & w7874) | (w7949 & w13420) | (w7874 & w13420);
assign w7974 = (~w7970 & w7973) | (~w7970 & w13037) | (w7973 & w13037);
assign w7975 = ~w7971 & ~w7974;
assign w7976 = A_442 & A_443;
assign w7977 = A_442 & ~A_443;
assign w7978 = ~A_442 & A_443;
assign w7979 = ~w7977 & ~w7978;
assign w7980 = (~w7976 & w7979) | (~w7976 & w12844) | (w7979 & w12844);
assign w7981 = A_439 & A_440;
assign w7982 = A_439 & ~A_440;
assign w7983 = ~A_439 & A_440;
assign w7984 = ~w7982 & ~w7983;
assign w7985 = (~w7981 & w7984) | (~w7981 & w12845) | (w7984 & w12845);
assign w7986 = w7980 & ~w7985;
assign w7987 = ~w7980 & w7985;
assign w7988 = A_441 & ~w7982;
assign w7989 = ~w7983 & w7988;
assign w7990 = ~A_441 & ~w7984;
assign w7991 = ~w7989 & ~w7990;
assign w7992 = A_444 & ~w7977;
assign w7993 = ~w7978 & w7992;
assign w7994 = ~A_444 & ~w7979;
assign w7995 = ~w7993 & ~w7994;
assign w7996 = ~w7991 & ~w7995;
assign w7997 = w7996 & w7998;
assign w7998 = ~w7986 & ~w7987;
assign w7999 = ~w7996 & ~w7998;
assign w8000 = ~w7997 & ~w7999;
assign w8001 = ~w7991 & w7995;
assign w8002 = w7991 & ~w7995;
assign w8003 = ~w8001 & ~w8002;
assign w8004 = w7996 & ~w7998;
assign w8005 = ~w7980 & ~w7985;
assign w8006 = ~w8004 & ~w8005;
assign w8007 = ~w8003 & ~w8006;
assign w8008 = ~w8000 & ~w8007;
assign w8009 = ~w8000 & ~w8006;
assign w8010 = A_448 & A_449;
assign w8011 = A_448 & ~A_449;
assign w8012 = ~A_448 & A_449;
assign w8013 = ~w8011 & ~w8012;
assign w8014 = (~w8010 & w8013) | (~w8010 & w12846) | (w8013 & w12846);
assign w8015 = A_445 & A_446;
assign w8016 = A_445 & ~A_446;
assign w8017 = ~A_445 & A_446;
assign w8018 = ~w8016 & ~w8017;
assign w8019 = (~w8015 & w8018) | (~w8015 & w12847) | (w8018 & w12847);
assign w8020 = ~w8014 & w8019;
assign w8021 = w8014 & ~w8019;
assign w8022 = ~w8020 & ~w8021;
assign w8023 = A_447 & ~w8016;
assign w8024 = ~w8017 & w8023;
assign w8025 = ~A_447 & ~w8018;
assign w8026 = ~w8024 & ~w8025;
assign w8027 = A_450 & ~w8011;
assign w8028 = ~w8012 & w8027;
assign w8029 = ~A_450 & ~w8013;
assign w8030 = ~w8028 & ~w8029;
assign w8031 = ~w8026 & ~w8030;
assign w8032 = ~w8022 & w8031;
assign w8033 = ~w8014 & ~w8019;
assign w8034 = ~w8032 & ~w8033;
assign w8035 = w8031 & w8022;
assign w8036 = ~w8022 & ~w8031;
assign w8037 = ~w8035 & ~w8036;
assign w8038 = ~w8034 & ~w8037;
assign w8039 = ~w8026 & w8030;
assign w8040 = w8026 & ~w8030;
assign w8041 = ~w8039 & ~w8040;
assign w8042 = ~w8003 & ~w8041;
assign w8043 = ~w8038 & w8042;
assign w8044 = ~w8009 & w8043;
assign w8045 = ~w8034 & ~w8041;
assign w8046 = ~w8037 & ~w8045;
assign w8047 = ~w8044 & w8046;
assign w8048 = w8044 & ~w8046;
assign w8049 = ~w8047 & ~w8048;
assign w8050 = ~w8008 & ~w8049;
assign w8051 = ~w8044 & ~w8046;
assign w8052 = ~w8037 & w8042;
assign w8053 = ~w8038 & w8052;
assign w8054 = ~w8009 & ~w8045;
assign w8055 = w8053 & w8054;
assign w8056 = (w8008 & w8051) | (w8008 & w13038) | (w8051 & w13038);
assign w8057 = ~w8050 & ~w8056;
assign w8058 = A_454 & A_455;
assign w8059 = A_454 & ~A_455;
assign w8060 = ~A_454 & A_455;
assign w8061 = ~w8059 & ~w8060;
assign w8062 = (~w8058 & w8061) | (~w8058 & w12848) | (w8061 & w12848);
assign w8063 = A_451 & A_452;
assign w8064 = A_451 & ~A_452;
assign w8065 = ~A_451 & A_452;
assign w8066 = ~w8064 & ~w8065;
assign w8067 = (~w8063 & w8066) | (~w8063 & w12849) | (w8066 & w12849);
assign w8068 = w8062 & ~w8067;
assign w8069 = ~w8062 & w8067;
assign w8070 = A_453 & ~w8064;
assign w8071 = ~w8065 & w8070;
assign w8072 = ~A_453 & ~w8066;
assign w8073 = ~w8071 & ~w8072;
assign w8074 = A_456 & ~w8059;
assign w8075 = ~w8060 & w8074;
assign w8076 = ~A_456 & ~w8061;
assign w8077 = ~w8075 & ~w8076;
assign w8078 = ~w8073 & ~w8077;
assign w8079 = w8078 & w8080;
assign w8080 = ~w8068 & ~w8069;
assign w8081 = ~w8078 & ~w8080;
assign w8082 = ~w8079 & ~w8081;
assign w8083 = ~w8073 & w8077;
assign w8084 = w8073 & ~w8077;
assign w8085 = ~w8083 & ~w8084;
assign w8086 = w8078 & ~w8080;
assign w8087 = ~w8062 & ~w8067;
assign w8088 = ~w8086 & ~w8087;
assign w8089 = ~w8085 & ~w8088;
assign w8090 = ~w8082 & ~w8089;
assign w8091 = ~w8082 & ~w8088;
assign w8092 = A_460 & A_461;
assign w8093 = A_460 & ~A_461;
assign w8094 = ~A_460 & A_461;
assign w8095 = ~w8093 & ~w8094;
assign w8096 = (~w8092 & w8095) | (~w8092 & w12850) | (w8095 & w12850);
assign w8097 = A_457 & A_458;
assign w8098 = A_457 & ~A_458;
assign w8099 = ~A_457 & A_458;
assign w8100 = ~w8098 & ~w8099;
assign w8101 = (~w8097 & w8100) | (~w8097 & w12851) | (w8100 & w12851);
assign w8102 = ~w8096 & w8101;
assign w8103 = w8096 & ~w8101;
assign w8104 = ~w8102 & ~w8103;
assign w8105 = A_459 & ~w8098;
assign w8106 = ~w8099 & w8105;
assign w8107 = ~A_459 & ~w8100;
assign w8108 = ~w8106 & ~w8107;
assign w8109 = A_462 & ~w8093;
assign w8110 = ~w8094 & w8109;
assign w8111 = ~A_462 & ~w8095;
assign w8112 = ~w8110 & ~w8111;
assign w8113 = ~w8108 & ~w8112;
assign w8114 = ~w8104 & w8113;
assign w8115 = ~w8096 & ~w8101;
assign w8116 = ~w8114 & ~w8115;
assign w8117 = w8113 & w8104;
assign w8118 = ~w8104 & ~w8113;
assign w8119 = ~w8117 & ~w8118;
assign w8120 = ~w8116 & ~w8119;
assign w8121 = ~w8108 & w8112;
assign w8122 = w8108 & ~w8112;
assign w8123 = ~w8121 & ~w8122;
assign w8124 = ~w8085 & ~w8123;
assign w8125 = ~w8120 & w8124;
assign w8126 = ~w8091 & w8125;
assign w8127 = ~w8116 & ~w8123;
assign w8128 = ~w8119 & ~w8127;
assign w8129 = ~w8126 & ~w8128;
assign w8130 = ~w8119 & w8124;
assign w8131 = ~w8120 & w8130;
assign w8132 = ~w8091 & ~w8127;
assign w8133 = w8131 & w8132;
assign w8134 = (w8090 & w8129) | (w8090 & w12852) | (w8129 & w12852);
assign w8135 = ~w8126 & w8128;
assign w8136 = w8126 & ~w8128;
assign w8137 = ~w8135 & ~w8136;
assign w8138 = ~w8090 & ~w8137;
assign w8139 = ~w8120 & ~w8123;
assign w8140 = ~w8085 & ~w8091;
assign w8141 = ~w8139 & w8140;
assign w8142 = w8139 & ~w8140;
assign w8143 = ~w8141 & ~w8142;
assign w8144 = ~w8038 & ~w8041;
assign w8145 = ~w8003 & ~w8009;
assign w8146 = ~w8144 & w8145;
assign w8147 = w8144 & ~w8145;
assign w8148 = ~w8146 & ~w8147;
assign w8149 = ~w8143 & ~w8148;
assign w8150 = ~w8138 & w12853;
assign w8151 = (w8149 & w8138) | (w8149 & w12854) | (w8138 & w12854);
assign w8152 = ~w8150 & ~w8151;
assign w8153 = ~w8057 & ~w8152;
assign w8154 = ~w8138 & w12855;
assign w8155 = (~w8149 & w8138) | (~w8149 & w13039) | (w8138 & w13039);
assign w8156 = (w8057 & w8155) | (w8057 & w12856) | (w8155 & w12856);
assign w8157 = ~w8143 & w8148;
assign w8158 = w8143 & ~w8148;
assign w8159 = ~w8157 & ~w8158;
assign w8160 = ~w7879 & w7948;
assign w8161 = w7879 & ~w7948;
assign w8162 = ~w8160 & ~w8161;
assign w8163 = ~w8159 & ~w8162;
assign w8164 = (~w12856 & w13040) | (~w12856 & w13041) | (w13040 & w13041);
assign w8165 = ~w8153 & w8164;
assign w8166 = ~w8153 & ~w8156;
assign w8167 = w8163 & ~w8166;
assign w8168 = (~w7975 & w8167) | (~w7975 & w13042) | (w8167 & w13042);
assign w8169 = w8163 & ~w8156;
assign w8170 = ~w8153 & w8169;
assign w8171 = ~w8163 & ~w8166;
assign w8172 = ~w8170 & ~w8171;
assign w8173 = (w7975 & w8171) | (w7975 & w13421) | (w8171 & w13421);
assign w8174 = ~w8159 & w8162;
assign w8175 = w8159 & ~w8162;
assign w8176 = ~w8174 & ~w8175;
assign w8177 = ~w7596 & w7737;
assign w8178 = w7596 & ~w7737;
assign w8179 = ~w8177 & ~w8178;
assign w8180 = ~w8176 & ~w8179;
assign w8181 = (~w8180 & w8172) | (~w8180 & w13043) | (w8172 & w13043);
assign w8182 = ~w8168 & w8181;
assign w8183 = (w8180 & w8173) | (w8180 & w13044) | (w8173 & w13044);
assign w8184 = ~w8182 & ~w8183;
assign w8185 = ~w7793 & ~w8184;
assign w8186 = (w8180 & w8172) | (w8180 & w13045) | (w8172 & w13045);
assign w8187 = ~w8168 & w8186;
assign w8188 = (~w8180 & w8173) | (~w8180 & w13046) | (w8173 & w13046);
assign w8189 = ~w8187 & ~w8188;
assign w8190 = w7793 & ~w8189;
assign w8191 = ~w8176 & w8179;
assign w8192 = w8176 & ~w8179;
assign w8193 = ~w8191 & ~w8192;
assign w8194 = ~w7016 & w7301;
assign w8195 = w7016 & ~w7301;
assign w8196 = ~w8194 & ~w8195;
assign w8197 = ~w8193 & ~w8196;
assign w8198 = (~w8197 & w8189) | (~w8197 & w13422) | (w8189 & w13422);
assign w8199 = ~w8185 & w8198;
assign w8200 = ~w8185 & ~w8190;
assign w8201 = w8197 & ~w8200;
assign w8202 = (~w7412 & w8201) | (~w7412 & w13423) | (w8201 & w13423);
assign w8203 = (w8197 & w8189) | (w8197 & w13881) | (w8189 & w13881);
assign w8204 = ~w8185 & w8203;
assign w8205 = ~w8197 & ~w8200;
assign w8206 = ~w8204 & ~w8205;
assign w8207 = (w7412 & w8205) | (w7412 & w13882) | (w8205 & w13882);
assign w8208 = ~w8193 & w8196;
assign w8209 = w8193 & ~w8196;
assign w8210 = ~w8208 & ~w8209;
assign w8211 = ~w5838 & w6411;
assign w8212 = w5838 & ~w6411;
assign w8213 = ~w8211 & ~w8212;
assign w8214 = ~w8210 & ~w8213;
assign w8215 = (~w8214 & w8206) | (~w8214 & w13424) | (w8206 & w13424);
assign w8216 = ~w8202 & w8215;
assign w8217 = (w8214 & w8207) | (w8214 & w13425) | (w8207 & w13425);
assign w8218 = ~w8216 & ~w8217;
assign w8219 = ~w6632 & ~w8218;
assign w8220 = (w8214 & w8206) | (w8214 & w13426) | (w8206 & w13426);
assign w8221 = ~w8202 & w8220;
assign w8222 = (~w8214 & w8207) | (~w8214 & w13427) | (w8207 & w13427);
assign w8223 = ~w8221 & ~w8222;
assign w8224 = w6632 & ~w8223;
assign w8225 = ~w8210 & w8213;
assign w8226 = w8210 & ~w8213;
assign w8227 = ~w8225 & ~w8226;
assign w8228 = ~w4262 & w4835;
assign w8229 = ~w4259 & ~w4835;
assign w8230 = ~w4261 & w8229;
assign w8231 = ~w8228 & ~w8230;
assign w8232 = ~w8227 & ~w8231;
assign w8233 = (~w8232 & w8223) | (~w8232 & w13883) | (w8223 & w13883);
assign w8234 = ~w8219 & w8233;
assign w8235 = ~w8219 & ~w8224;
assign w8236 = w8232 & ~w8235;
assign w8237 = (~w5056 & w8236) | (~w5056 & w13884) | (w8236 & w13884);
assign w8238 = ~w2720 & w2723;
assign w8239 = w2720 & ~w2723;
assign w8240 = ~w8238 & ~w8239;
assign w8241 = ~w8227 & w8231;
assign w8242 = w8227 & ~w8231;
assign w8243 = ~w8241 & ~w8242;
assign w8244 = ~w8240 & ~w8243;
assign w8245 = (w8232 & w8223) | (w8232 & w13885) | (w8223 & w13885);
assign w8246 = ~w8219 & w8245;
assign w8247 = ~w8232 & ~w8235;
assign w8248 = (w5056 & w8247) | (w5056 & w13886) | (w8247 & w13886);
assign w8249 = ~w8244 & ~w8248;
assign w8250 = ~w8237 & w8249;
assign w8251 = (~w3162 & ~w8249) | (~w3162 & w13887) | (~w8249 & w13887);
assign w8252 = ~w8237 & ~w8248;
assign w8253 = w8244 & ~w8252;
assign w8254 = ~w8251 & ~w8253;
assign w8255 = ~w5056 & ~w8234;
assign w8256 = ~w8236 & ~w8255;
assign w8257 = (~w5049 & ~w5051) | (~w5049 & w12857) | (~w5051 & w12857);
assign w8258 = ~w5053 & ~w8257;
assign w8259 = (~w3542 & ~w4249) | (~w3542 & w12858) | (~w4249 & w12858);
assign w8260 = ~w4252 & ~w8259;
assign w8261 = ~w3842 & ~w4233;
assign w8262 = ~w4234 & ~w8261;
assign w8263 = ~w3836 & ~w3839;
assign w8264 = ~w3840 & ~w8263;
assign w8265 = (w3801 & ~w3831) | (w3801 & w12859) | (~w3831 & w12859);
assign w8266 = ~w3833 & ~w8265;
assign w8267 = (~w3818 & w3814) | (~w3818 & w12860) | (w3814 & w12860);
assign w8268 = ~w3816 & ~w8267;
assign w8269 = ~w3805 & ~w3807;
assign w8270 = ~w3813 & ~w8269;
assign w8271 = ~w8268 & w8270;
assign w8272 = ~w3816 & ~w8270;
assign w8273 = ~w8267 & w8272;
assign w8274 = ~w3743 & ~w3757;
assign w8275 = ~w3754 & ~w8274;
assign w8276 = (w8275 & ~w8272) | (w8275 & w12861) | (~w8272 & w12861);
assign w8277 = ~w8271 & w8276;
assign w8278 = ~w8271 & ~w8273;
assign w8279 = ~w8275 & ~w8278;
assign w8280 = ~w8277 & ~w8279;
assign w8281 = ~w8266 & ~w8280;
assign w8282 = ~w3833 & ~w8277;
assign w8283 = w8282 & w12862;
assign w8284 = ~w8281 & ~w8283;
assign w8285 = ~w3624 & ~w3717;
assign w8286 = ~w3718 & ~w8285;
assign w8287 = (w3575 & w3611) | (w3575 & w13047) | (w3611 & w13047);
assign w8288 = ~w3622 & ~w8287;
assign w8289 = ~w3604 & ~w3608;
assign w8290 = ~w3601 & ~w8289;
assign w8291 = ~w3567 & ~w3570;
assign w8292 = ~w3573 & ~w8291;
assign w8293 = ~w8290 & w8292;
assign w8294 = w8290 & ~w8292;
assign w8295 = ~w8293 & ~w8294;
assign w8296 = ~w8288 & ~w8295;
assign w8297 = ~w3622 & ~w8293;
assign w8298 = ~w8294 & w8297;
assign w8299 = ~w8287 & w8298;
assign w8300 = ~w8296 & ~w8299;
assign w8301 = (w3657 & w3693) | (w3657 & w13048) | (w3693 & w13048);
assign w8302 = ~w3700 & ~w8301;
assign w8303 = ~w3686 & ~w3690;
assign w8304 = ~w3683 & ~w8303;
assign w8305 = ~w3649 & ~w3652;
assign w8306 = ~w3655 & ~w8305;
assign w8307 = ~w8304 & w8306;
assign w8308 = w8304 & ~w8306;
assign w8309 = ~w8307 & ~w8308;
assign w8310 = ~w8302 & ~w8309;
assign w8311 = ~w3700 & ~w8307;
assign w8312 = ~w8308 & w8311;
assign w8313 = ~w8301 & w8312;
assign w8314 = ~w8310 & ~w8313;
assign w8315 = ~w8300 & w8314;
assign w8316 = w8300 & ~w8314;
assign w8317 = ~w8315 & ~w8316;
assign w8318 = ~w8286 & ~w8317;
assign w8319 = w8286 & w8317;
assign w8320 = ~w8318 & ~w8319;
assign w8321 = ~w8284 & w8320;
assign w8322 = w8284 & ~w8320;
assign w8323 = ~w8321 & ~w8322;
assign w8324 = ~w8264 & ~w8323;
assign w8325 = w8264 & w8323;
assign w8326 = ~w8324 & ~w8325;
assign w8327 = ~w4025 & ~w4215;
assign w8328 = ~w4217 & ~w8327;
assign w8329 = ~w4019 & ~w4021;
assign w8330 = ~w4022 & ~w8329;
assign w8331 = (w4003 & w4006) | (w4003 & w12863) | (w4006 & w12863);
assign w8332 = ~w4017 & ~w8331;
assign w8333 = ~w3945 & ~w3959;
assign w8334 = ~w3956 & ~w8333;
assign w8335 = ~w3978 & ~w3992;
assign w8336 = ~w3989 & ~w8335;
assign w8337 = ~w8334 & w8336;
assign w8338 = w8334 & ~w8336;
assign w8339 = ~w8337 & ~w8338;
assign w8340 = ~w8332 & ~w8339;
assign w8341 = ~w4017 & ~w8337;
assign w8342 = ~w8338 & w8341;
assign w8343 = ~w8331 & w8342;
assign w8344 = ~w8340 & ~w8343;
assign w8345 = (w3875 & w3911) | (w3875 & w12864) | (w3911 & w12864);
assign w8346 = ~w3918 & ~w8345;
assign w8347 = ~w3904 & ~w3908;
assign w8348 = ~w3901 & ~w8347;
assign w8349 = ~w3867 & ~w3870;
assign w8350 = ~w3873 & ~w8349;
assign w8351 = ~w8348 & w8350;
assign w8352 = w8348 & ~w8350;
assign w8353 = ~w8351 & ~w8352;
assign w8354 = ~w8346 & ~w8353;
assign w8355 = ~w3918 & ~w8351;
assign w8356 = ~w8352 & w8355;
assign w8357 = ~w8345 & w8356;
assign w8358 = ~w8354 & ~w8357;
assign w8359 = ~w8344 & w8358;
assign w8360 = w8344 & ~w8358;
assign w8361 = ~w8359 & ~w8360;
assign w8362 = ~w8330 & ~w8361;
assign w8363 = w8330 & w8361;
assign w8364 = ~w8362 & ~w8363;
assign w8365 = ~w4107 & ~w4200;
assign w8366 = ~w4201 & ~w8365;
assign w8367 = (w4058 & w4094) | (w4058 & w12865) | (w4094 & w12865);
assign w8368 = ~w4105 & ~w8367;
assign w8369 = ~w4087 & ~w4091;
assign w8370 = ~w4084 & ~w8369;
assign w8371 = ~w4050 & ~w4053;
assign w8372 = ~w4056 & ~w8371;
assign w8373 = ~w8370 & w8372;
assign w8374 = w8370 & ~w8372;
assign w8375 = ~w8373 & ~w8374;
assign w8376 = ~w8368 & ~w8375;
assign w8377 = ~w4105 & ~w8373;
assign w8378 = ~w8374 & w8377;
assign w8379 = ~w8367 & w8378;
assign w8380 = ~w8376 & ~w8379;
assign w8381 = (w4140 & w4176) | (w4140 & w12866) | (w4176 & w12866);
assign w8382 = ~w4183 & ~w8381;
assign w8383 = ~w4169 & ~w4173;
assign w8384 = ~w4166 & ~w8383;
assign w8385 = ~w4132 & ~w4135;
assign w8386 = ~w4138 & ~w8385;
assign w8387 = ~w8384 & w8386;
assign w8388 = w8384 & ~w8386;
assign w8389 = ~w8387 & ~w8388;
assign w8390 = ~w8382 & ~w8389;
assign w8391 = ~w4183 & ~w8387;
assign w8392 = ~w8388 & w8391;
assign w8393 = ~w8381 & w8392;
assign w8394 = ~w8390 & ~w8393;
assign w8395 = ~w8380 & w8394;
assign w8396 = w8380 & ~w8394;
assign w8397 = ~w8395 & ~w8396;
assign w8398 = ~w8366 & ~w8397;
assign w8399 = w8366 & w8397;
assign w8400 = ~w8398 & ~w8399;
assign w8401 = ~w8364 & w8400;
assign w8402 = w8364 & ~w8400;
assign w8403 = ~w8401 & ~w8402;
assign w8404 = ~w8328 & ~w8403;
assign w8405 = w8328 & w8403;
assign w8406 = ~w8404 & ~w8405;
assign w8407 = ~w8326 & w8406;
assign w8408 = w8326 & ~w8406;
assign w8409 = ~w8407 & ~w8408;
assign w8410 = w8262 & w8409;
assign w8411 = ~w8262 & ~w8409;
assign w8412 = ~w3536 & ~w3539;
assign w8413 = ~w3540 & ~w8412;
assign w8414 = ~w3531 & ~w3533;
assign w8415 = ~w3534 & ~w8414;
assign w8416 = (w3515 & w3518) | (w3515 & w13733) | (w3518 & w13733);
assign w8417 = ~w3529 & ~w8416;
assign w8418 = ~w3432 & ~w3446;
assign w8419 = ~w3443 & ~w8418;
assign w8420 = ~w3465 & ~w3479;
assign w8421 = ~w3476 & ~w8420;
assign w8422 = ~w8419 & w8421;
assign w8423 = w8419 & ~w8421;
assign w8424 = ~w8422 & ~w8423;
assign w8425 = ~w8417 & ~w8424;
assign w8426 = ~w3529 & ~w8422;
assign w8427 = ~w8423 & w8426;
assign w8428 = ~w8416 & w8427;
assign w8429 = ~w8425 & ~w8428;
assign w8430 = (w3494 & w3497) | (w3494 & w13734) | (w3497 & w13734);
assign w8431 = ~w3504 & ~w8430;
assign w8432 = ~w3363 & ~w3377;
assign w8433 = ~w3374 & ~w8432;
assign w8434 = ~w3396 & ~w3410;
assign w8435 = ~w3407 & ~w8434;
assign w8436 = ~w8433 & w8435;
assign w8437 = w8433 & ~w8435;
assign w8438 = ~w8436 & ~w8437;
assign w8439 = ~w8431 & ~w8438;
assign w8440 = ~w3504 & ~w8436;
assign w8441 = ~w8437 & w8440;
assign w8442 = ~w8430 & w8441;
assign w8443 = ~w8439 & ~w8442;
assign w8444 = ~w8429 & w8443;
assign w8445 = w8429 & ~w8443;
assign w8446 = ~w8444 & ~w8445;
assign w8447 = ~w8415 & ~w8446;
assign w8448 = w8415 & w8446;
assign w8449 = ~w8447 & ~w8448;
assign w8450 = ~w3244 & ~w3337;
assign w8451 = ~w3338 & ~w8450;
assign w8452 = (w3195 & w3231) | (w3195 & w13735) | (w3231 & w13735);
assign w8453 = ~w3242 & ~w8452;
assign w8454 = ~w3224 & ~w3228;
assign w8455 = ~w3221 & ~w8454;
assign w8456 = ~w3187 & ~w3190;
assign w8457 = ~w3193 & ~w8456;
assign w8458 = ~w8455 & w8457;
assign w8459 = w8455 & ~w8457;
assign w8460 = ~w8458 & ~w8459;
assign w8461 = ~w8453 & ~w8460;
assign w8462 = ~w3242 & ~w8458;
assign w8463 = ~w8459 & w8462;
assign w8464 = ~w8452 & w8463;
assign w8465 = ~w8461 & ~w8464;
assign w8466 = (w3277 & w3313) | (w3277 & w13736) | (w3313 & w13736);
assign w8467 = ~w3320 & ~w8466;
assign w8468 = ~w3306 & ~w3310;
assign w8469 = ~w3303 & ~w8468;
assign w8470 = ~w3269 & ~w3272;
assign w8471 = ~w3275 & ~w8470;
assign w8472 = ~w8469 & w8471;
assign w8473 = w8469 & ~w8471;
assign w8474 = ~w8472 & ~w8473;
assign w8475 = ~w8467 & ~w8474;
assign w8476 = ~w3320 & ~w8472;
assign w8477 = ~w8473 & w8476;
assign w8478 = ~w8466 & w8477;
assign w8479 = ~w8475 & ~w8478;
assign w8480 = ~w8465 & w8479;
assign w8481 = w8465 & ~w8479;
assign w8482 = ~w8480 & ~w8481;
assign w8483 = ~w8451 & ~w8482;
assign w8484 = w8451 & w8482;
assign w8485 = ~w8483 & ~w8484;
assign w8486 = ~w8449 & w8485;
assign w8487 = w8449 & ~w8485;
assign w8488 = ~w8486 & ~w8487;
assign w8489 = ~w8413 & ~w8488;
assign w8490 = w8413 & w8488;
assign w8491 = ~w8489 & ~w8490;
assign w8492 = (~w8491 & w8409) | (~w8491 & w13539) | (w8409 & w13539);
assign w8493 = ~w8410 & w8492;
assign w8494 = ~w8410 & ~w8411;
assign w8495 = w8491 & ~w8494;
assign w8496 = ~w8493 & ~w8495;
assign w8497 = ~w8495 & w13540;
assign w8498 = (~w8260 & w8495) | (~w8260 & w13541) | (w8495 & w13541);
assign w8499 = ~w5042 & ~w5045;
assign w8500 = ~w5046 & ~w8499;
assign w8501 = ~w5036 & ~w5039;
assign w8502 = ~w5040 & ~w8501;
assign w8503 = ~w5031 & ~w5033;
assign w8504 = ~w5034 & ~w8503;
assign w8505 = (w5015 & w5018) | (w5015 & w13542) | (w5018 & w13542);
assign w8506 = ~w5029 & ~w8505;
assign w8507 = ~w4774 & ~w4788;
assign w8508 = ~w4785 & ~w8507;
assign w8509 = ~w4807 & ~w4821;
assign w8510 = ~w4818 & ~w8509;
assign w8511 = ~w8508 & w8510;
assign w8512 = w8508 & ~w8510;
assign w8513 = ~w8511 & ~w8512;
assign w8514 = ~w8506 & ~w8513;
assign w8515 = ~w5029 & ~w8511;
assign w8516 = ~w8512 & w8515;
assign w8517 = ~w8505 & w8516;
assign w8518 = ~w8514 & ~w8517;
assign w8519 = (w4994 & w4997) | (w4994 & w13543) | (w4997 & w13543);
assign w8520 = ~w5004 & ~w8519;
assign w8521 = ~w4705 & ~w4719;
assign w8522 = ~w4716 & ~w8521;
assign w8523 = ~w4738 & ~w4752;
assign w8524 = ~w4749 & ~w8523;
assign w8525 = ~w8522 & w8524;
assign w8526 = w8522 & ~w8524;
assign w8527 = ~w8525 & ~w8526;
assign w8528 = ~w8520 & ~w8527;
assign w8529 = ~w5004 & ~w8525;
assign w8530 = ~w8526 & w8529;
assign w8531 = ~w8519 & w8530;
assign w8532 = ~w8528 & ~w8531;
assign w8533 = ~w8518 & w8532;
assign w8534 = w8518 & ~w8532;
assign w8535 = ~w8533 & ~w8534;
assign w8536 = ~w8504 & ~w8535;
assign w8537 = w8504 & w8535;
assign w8538 = ~w8536 & ~w8537;
assign w8539 = ~w4962 & ~w4981;
assign w8540 = ~w4982 & ~w8539;
assign w8541 = (w4946 & w4949) | (w4946 & w13544) | (w4949 & w13544);
assign w8542 = ~w4960 & ~w8541;
assign w8543 = ~w4633 & ~w4647;
assign w8544 = ~w4644 & ~w8543;
assign w8545 = ~w4666 & ~w4680;
assign w8546 = ~w4677 & ~w8545;
assign w8547 = ~w8544 & w8546;
assign w8548 = w8544 & ~w8546;
assign w8549 = ~w8547 & ~w8548;
assign w8550 = ~w8542 & ~w8549;
assign w8551 = ~w4960 & ~w8547;
assign w8552 = ~w8548 & w8551;
assign w8553 = ~w8541 & w8552;
assign w8554 = ~w8550 & ~w8553;
assign w8555 = (w4964 & w4967) | (w4964 & w13545) | (w4967 & w13545);
assign w8556 = ~w4974 & ~w8555;
assign w8557 = ~w4564 & ~w4578;
assign w8558 = ~w4575 & ~w8557;
assign w8559 = ~w4597 & ~w4611;
assign w8560 = ~w4608 & ~w8559;
assign w8561 = ~w8558 & w8560;
assign w8562 = w8558 & ~w8560;
assign w8563 = ~w8561 & ~w8562;
assign w8564 = ~w8556 & ~w8563;
assign w8565 = ~w4974 & ~w8561;
assign w8566 = ~w8562 & w8565;
assign w8567 = ~w8555 & w8566;
assign w8568 = ~w8564 & ~w8567;
assign w8569 = ~w8554 & w8568;
assign w8570 = w8554 & ~w8568;
assign w8571 = ~w8569 & ~w8570;
assign w8572 = ~w8540 & ~w8571;
assign w8573 = w8540 & w8571;
assign w8574 = ~w8572 & ~w8573;
assign w8575 = ~w8538 & w8574;
assign w8576 = w8538 & ~w8574;
assign w8577 = ~w8575 & ~w8576;
assign w8578 = ~w8502 & ~w8577;
assign w8579 = w8502 & w8577;
assign w8580 = ~w8578 & ~w8579;
assign w8581 = ~w4885 & ~w4931;
assign w8582 = ~w4933 & ~w8581;
assign w8583 = ~w4880 & ~w4882;
assign w8584 = ~w4883 & ~w8583;
assign w8585 = (w4864 & w4867) | (w4864 & w13546) | (w4867 & w13546);
assign w8586 = ~w4878 & ~w8585;
assign w8587 = ~w4489 & ~w4503;
assign w8588 = ~w4500 & ~w8587;
assign w8589 = ~w4522 & ~w4536;
assign w8590 = ~w4533 & ~w8589;
assign w8591 = ~w8588 & w8590;
assign w8592 = w8588 & ~w8590;
assign w8593 = ~w8591 & ~w8592;
assign w8594 = ~w8586 & ~w8593;
assign w8595 = ~w4878 & ~w8591;
assign w8596 = ~w8592 & w8595;
assign w8597 = ~w8585 & w8596;
assign w8598 = ~w8594 & ~w8597;
assign w8599 = (w4843 & w4846) | (w4843 & w13547) | (w4846 & w13547);
assign w8600 = ~w4853 & ~w8599;
assign w8601 = ~w4420 & ~w4434;
assign w8602 = ~w4431 & ~w8601;
assign w8603 = ~w4453 & ~w4467;
assign w8604 = ~w4464 & ~w8603;
assign w8605 = ~w8602 & w8604;
assign w8606 = w8602 & ~w8604;
assign w8607 = ~w8605 & ~w8606;
assign w8608 = ~w8600 & ~w8607;
assign w8609 = ~w4853 & ~w8605;
assign w8610 = ~w8606 & w8609;
assign w8611 = ~w8599 & w8610;
assign w8612 = ~w8608 & ~w8611;
assign w8613 = ~w8598 & w8612;
assign w8614 = w8598 & ~w8612;
assign w8615 = ~w8613 & ~w8614;
assign w8616 = ~w8584 & ~w8615;
assign w8617 = w8584 & w8615;
assign w8618 = ~w8616 & ~w8617;
assign w8619 = ~w4903 & ~w4922;
assign w8620 = ~w4923 & ~w8619;
assign w8621 = (w4887 & w4890) | (w4887 & w13548) | (w4890 & w13548);
assign w8622 = ~w4901 & ~w8621;
assign w8623 = ~w4348 & ~w4362;
assign w8624 = ~w4359 & ~w8623;
assign w8625 = ~w4381 & ~w4395;
assign w8626 = ~w4392 & ~w8625;
assign w8627 = ~w8624 & w8626;
assign w8628 = w8624 & ~w8626;
assign w8629 = ~w8627 & ~w8628;
assign w8630 = ~w8622 & ~w8629;
assign w8631 = ~w4901 & ~w8627;
assign w8632 = ~w8628 & w8631;
assign w8633 = ~w8621 & w8632;
assign w8634 = ~w8630 & ~w8633;
assign w8635 = (w4905 & w4908) | (w4905 & w13549) | (w4908 & w13549);
assign w8636 = ~w4915 & ~w8635;
assign w8637 = ~w4279 & ~w4293;
assign w8638 = ~w4290 & ~w8637;
assign w8639 = ~w4312 & ~w4326;
assign w8640 = ~w4323 & ~w8639;
assign w8641 = ~w8638 & w8640;
assign w8642 = w8638 & ~w8640;
assign w8643 = ~w8641 & ~w8642;
assign w8644 = ~w8636 & ~w8643;
assign w8645 = ~w4915 & ~w8641;
assign w8646 = ~w8642 & w8645;
assign w8647 = ~w8635 & w8646;
assign w8648 = ~w8644 & ~w8647;
assign w8649 = ~w8634 & w8648;
assign w8650 = w8634 & ~w8648;
assign w8651 = ~w8649 & ~w8650;
assign w8652 = ~w8620 & ~w8651;
assign w8653 = w8620 & w8651;
assign w8654 = ~w8652 & ~w8653;
assign w8655 = ~w8618 & w8654;
assign w8656 = w8618 & ~w8654;
assign w8657 = ~w8655 & ~w8656;
assign w8658 = ~w8582 & ~w8657;
assign w8659 = w8582 & w8657;
assign w8660 = ~w8658 & ~w8659;
assign w8661 = ~w8580 & w8660;
assign w8662 = w8580 & ~w8660;
assign w8663 = ~w8661 & ~w8662;
assign w8664 = ~w8500 & ~w8663;
assign w8665 = w8500 & w8663;
assign w8666 = ~w8664 & ~w8665;
assign w8667 = (~w8666 & w8496) | (~w8666 & w12867) | (w8496 & w12867);
assign w8668 = ~w8497 & w8667;
assign w8669 = ~w8497 & ~w8498;
assign w8670 = w8666 & ~w8669;
assign w8671 = (~w8258 & w8670) | (~w8258 & w13428) | (w8670 & w13428);
assign w8672 = ~w8670 & w13429;
assign w8673 = ~w8671 & ~w8672;
assign w8674 = ~w6632 & ~w8216;
assign w8675 = ~w8217 & ~w8674;
assign w8676 = ~w6626 & ~w6629;
assign w8677 = ~w6630 & ~w8676;
assign w8678 = ~w6619 & ~w6622;
assign w8679 = ~w6623 & ~w8678;
assign w8680 = ~w6613 & ~w6616;
assign w8681 = ~w6617 & ~w8680;
assign w8682 = ~w6607 & ~w6609;
assign w8683 = ~w6610 & ~w8682;
assign w8684 = (w6591 & w6594) | (w6591 & w12868) | (w6594 & w12868);
assign w8685 = ~w6605 & ~w8684;
assign w8686 = ~w6350 & ~w6364;
assign w8687 = ~w6361 & ~w8686;
assign w8688 = ~w6383 & ~w6397;
assign w8689 = ~w6394 & ~w8688;
assign w8690 = ~w8687 & w8689;
assign w8691 = w8687 & ~w8689;
assign w8692 = ~w8690 & ~w8691;
assign w8693 = ~w8685 & ~w8692;
assign w8694 = ~w6605 & ~w8690;
assign w8695 = ~w8691 & w8694;
assign w8696 = ~w8684 & w8695;
assign w8697 = ~w8693 & ~w8696;
assign w8698 = (w6570 & w6573) | (w6570 & w12869) | (w6573 & w12869);
assign w8699 = ~w6580 & ~w8698;
assign w8700 = ~w6281 & ~w6295;
assign w8701 = ~w6292 & ~w8700;
assign w8702 = ~w6314 & ~w6328;
assign w8703 = ~w6325 & ~w8702;
assign w8704 = ~w8701 & w8703;
assign w8705 = w8701 & ~w8703;
assign w8706 = ~w8704 & ~w8705;
assign w8707 = ~w8699 & ~w8706;
assign w8708 = ~w6580 & ~w8704;
assign w8709 = ~w8705 & w8708;
assign w8710 = ~w8698 & w8709;
assign w8711 = ~w8707 & ~w8710;
assign w8712 = ~w8697 & w8711;
assign w8713 = w8697 & ~w8711;
assign w8714 = ~w8712 & ~w8713;
assign w8715 = ~w8683 & ~w8714;
assign w8716 = w8683 & w8714;
assign w8717 = ~w8715 & ~w8716;
assign w8718 = ~w6538 & ~w6557;
assign w8719 = ~w6558 & ~w8718;
assign w8720 = (w6522 & w6525) | (w6522 & w12870) | (w6525 & w12870);
assign w8721 = ~w6536 & ~w8720;
assign w8722 = ~w6209 & ~w6223;
assign w8723 = ~w6220 & ~w8722;
assign w8724 = ~w6242 & ~w6256;
assign w8725 = ~w6253 & ~w8724;
assign w8726 = ~w8723 & w8725;
assign w8727 = w8723 & ~w8725;
assign w8728 = ~w8726 & ~w8727;
assign w8729 = ~w8721 & ~w8728;
assign w8730 = ~w6536 & ~w8726;
assign w8731 = ~w8727 & w8730;
assign w8732 = ~w8720 & w8731;
assign w8733 = ~w8729 & ~w8732;
assign w8734 = (w6540 & w6543) | (w6540 & w12871) | (w6543 & w12871);
assign w8735 = ~w6550 & ~w8734;
assign w8736 = ~w6140 & ~w6154;
assign w8737 = ~w6151 & ~w8736;
assign w8738 = ~w6173 & ~w6187;
assign w8739 = ~w6184 & ~w8738;
assign w8740 = ~w8737 & w8739;
assign w8741 = w8737 & ~w8739;
assign w8742 = ~w8740 & ~w8741;
assign w8743 = ~w8735 & ~w8742;
assign w8744 = ~w6550 & ~w8740;
assign w8745 = ~w8741 & w8744;
assign w8746 = ~w8734 & w8745;
assign w8747 = ~w8743 & ~w8746;
assign w8748 = ~w8733 & w8747;
assign w8749 = w8733 & ~w8747;
assign w8750 = ~w8748 & ~w8749;
assign w8751 = ~w8719 & ~w8750;
assign w8752 = w8719 & w8750;
assign w8753 = ~w8751 & ~w8752;
assign w8754 = ~w8717 & w8753;
assign w8755 = w8717 & ~w8753;
assign w8756 = ~w8754 & ~w8755;
assign w8757 = ~w8681 & ~w8756;
assign w8758 = w8681 & w8756;
assign w8759 = ~w8757 & ~w8758;
assign w8760 = ~w6461 & ~w6507;
assign w8761 = ~w6509 & ~w8760;
assign w8762 = ~w6455 & ~w6457;
assign w8763 = ~w6458 & ~w8762;
assign w8764 = (w6439 & w6442) | (w6439 & w12872) | (w6442 & w12872);
assign w8765 = ~w6453 & ~w8764;
assign w8766 = ~w6065 & ~w6079;
assign w8767 = ~w6076 & ~w8766;
assign w8768 = ~w6098 & ~w6112;
assign w8769 = ~w6109 & ~w8768;
assign w8770 = ~w8767 & w8769;
assign w8771 = w8767 & ~w8769;
assign w8772 = ~w8770 & ~w8771;
assign w8773 = ~w8765 & ~w8772;
assign w8774 = ~w6453 & ~w8770;
assign w8775 = ~w8771 & w8774;
assign w8776 = ~w8764 & w8775;
assign w8777 = ~w8773 & ~w8776;
assign w8778 = (w6418 & w6421) | (w6418 & w12873) | (w6421 & w12873);
assign w8779 = ~w6428 & ~w8778;
assign w8780 = ~w5996 & ~w6010;
assign w8781 = ~w6007 & ~w8780;
assign w8782 = ~w6029 & ~w6043;
assign w8783 = ~w6040 & ~w8782;
assign w8784 = ~w8781 & w8783;
assign w8785 = w8781 & ~w8783;
assign w8786 = ~w8784 & ~w8785;
assign w8787 = ~w8779 & ~w8786;
assign w8788 = ~w6428 & ~w8784;
assign w8789 = ~w8785 & w8788;
assign w8790 = ~w8778 & w8789;
assign w8791 = ~w8787 & ~w8790;
assign w8792 = ~w8777 & w8791;
assign w8793 = w8777 & ~w8791;
assign w8794 = ~w8792 & ~w8793;
assign w8795 = ~w8763 & ~w8794;
assign w8796 = w8763 & w8794;
assign w8797 = ~w8795 & ~w8796;
assign w8798 = ~w6479 & ~w6498;
assign w8799 = ~w6499 & ~w8798;
assign w8800 = (w6463 & w6466) | (w6463 & w12874) | (w6466 & w12874);
assign w8801 = ~w6477 & ~w8800;
assign w8802 = ~w5924 & ~w5938;
assign w8803 = ~w5935 & ~w8802;
assign w8804 = ~w5957 & ~w5971;
assign w8805 = ~w5968 & ~w8804;
assign w8806 = ~w8803 & w8805;
assign w8807 = w8803 & ~w8805;
assign w8808 = ~w8806 & ~w8807;
assign w8809 = ~w8801 & ~w8808;
assign w8810 = ~w6477 & ~w8806;
assign w8811 = ~w8807 & w8810;
assign w8812 = ~w8800 & w8811;
assign w8813 = ~w8809 & ~w8812;
assign w8814 = (w6481 & w6484) | (w6481 & w12875) | (w6484 & w12875);
assign w8815 = ~w6491 & ~w8814;
assign w8816 = ~w5855 & ~w5869;
assign w8817 = ~w5866 & ~w8816;
assign w8818 = ~w5888 & ~w5902;
assign w8819 = ~w5899 & ~w8818;
assign w8820 = ~w8817 & w8819;
assign w8821 = w8817 & ~w8819;
assign w8822 = ~w8820 & ~w8821;
assign w8823 = ~w8815 & ~w8822;
assign w8824 = ~w6491 & ~w8820;
assign w8825 = ~w8821 & w8824;
assign w8826 = ~w8814 & w8825;
assign w8827 = ~w8823 & ~w8826;
assign w8828 = ~w8813 & w8827;
assign w8829 = w8813 & ~w8827;
assign w8830 = ~w8828 & ~w8829;
assign w8831 = ~w8799 & ~w8830;
assign w8832 = w8799 & w8830;
assign w8833 = ~w8831 & ~w8832;
assign w8834 = ~w8797 & w8833;
assign w8835 = w8797 & ~w8833;
assign w8836 = ~w8834 & ~w8835;
assign w8837 = ~w8761 & ~w8836;
assign w8838 = w8761 & w8836;
assign w8839 = ~w8837 & ~w8838;
assign w8840 = ~w8759 & w8839;
assign w8841 = w8759 & ~w8839;
assign w8842 = ~w8840 & ~w8841;
assign w8843 = ~w8679 & ~w8842;
assign w8844 = w8679 & w8842;
assign w8845 = ~w8843 & ~w8844;
assign w8846 = ~w5437 & ~w5827;
assign w8847 = ~w5828 & ~w8846;
assign w8848 = ~w5431 & ~w5434;
assign w8849 = ~w5435 & ~w8848;
assign w8850 = ~w5425 & ~w5427;
assign w8851 = ~w5428 & ~w8850;
assign w8852 = (w5409 & w5412) | (w5409 & w12876) | (w5412 & w12876);
assign w8853 = ~w5423 & ~w8852;
assign w8854 = ~w5326 & ~w5340;
assign w8855 = ~w5337 & ~w8854;
assign w8856 = ~w5359 & ~w5373;
assign w8857 = ~w5370 & ~w8856;
assign w8858 = ~w8855 & w8857;
assign w8859 = w8855 & ~w8857;
assign w8860 = ~w8858 & ~w8859;
assign w8861 = ~w8853 & ~w8860;
assign w8862 = ~w5423 & ~w8858;
assign w8863 = ~w8859 & w8862;
assign w8864 = ~w8852 & w8863;
assign w8865 = ~w8861 & ~w8864;
assign w8866 = (w5388 & w5391) | (w5388 & w12877) | (w5391 & w12877);
assign w8867 = ~w5398 & ~w8866;
assign w8868 = ~w5257 & ~w5271;
assign w8869 = ~w5268 & ~w8868;
assign w8870 = ~w5290 & ~w5304;
assign w8871 = ~w5301 & ~w8870;
assign w8872 = ~w8869 & w8871;
assign w8873 = w8869 & ~w8871;
assign w8874 = ~w8872 & ~w8873;
assign w8875 = ~w8867 & ~w8874;
assign w8876 = ~w5398 & ~w8872;
assign w8877 = ~w8873 & w8876;
assign w8878 = ~w8866 & w8877;
assign w8879 = ~w8875 & ~w8878;
assign w8880 = ~w8865 & w8879;
assign w8881 = w8865 & ~w8879;
assign w8882 = ~w8880 & ~w8881;
assign w8883 = ~w8851 & ~w8882;
assign w8884 = w8851 & w8882;
assign w8885 = ~w8883 & ~w8884;
assign w8886 = ~w5138 & ~w5231;
assign w8887 = ~w5232 & ~w8886;
assign w8888 = (w5089 & w5125) | (w5089 & w12878) | (w5125 & w12878);
assign w8889 = ~w5136 & ~w8888;
assign w8890 = ~w5118 & ~w5122;
assign w8891 = ~w5115 & ~w8890;
assign w8892 = ~w5081 & ~w5084;
assign w8893 = ~w5087 & ~w8892;
assign w8894 = ~w8891 & w8893;
assign w8895 = w8891 & ~w8893;
assign w8896 = ~w8894 & ~w8895;
assign w8897 = ~w8889 & ~w8896;
assign w8898 = ~w5136 & ~w8894;
assign w8899 = ~w8895 & w8898;
assign w8900 = ~w8888 & w8899;
assign w8901 = ~w8897 & ~w8900;
assign w8902 = (w5171 & w5207) | (w5171 & w12879) | (w5207 & w12879);
assign w8903 = ~w5214 & ~w8902;
assign w8904 = ~w5200 & ~w5204;
assign w8905 = ~w5197 & ~w8904;
assign w8906 = ~w5163 & ~w5166;
assign w8907 = ~w5169 & ~w8906;
assign w8908 = ~w8905 & w8907;
assign w8909 = w8905 & ~w8907;
assign w8910 = ~w8908 & ~w8909;
assign w8911 = ~w8903 & ~w8910;
assign w8912 = ~w5214 & ~w8908;
assign w8913 = ~w8909 & w8912;
assign w8914 = ~w8902 & w8913;
assign w8915 = ~w8911 & ~w8914;
assign w8916 = ~w8901 & w8915;
assign w8917 = w8901 & ~w8915;
assign w8918 = ~w8916 & ~w8917;
assign w8919 = ~w8887 & ~w8918;
assign w8920 = w8887 & w8918;
assign w8921 = ~w8919 & ~w8920;
assign w8922 = ~w8885 & w8921;
assign w8923 = w8885 & ~w8921;
assign w8924 = ~w8922 & ~w8923;
assign w8925 = ~w8849 & ~w8924;
assign w8926 = w8849 & w8924;
assign w8927 = ~w8925 & ~w8926;
assign w8928 = ~w5620 & ~w5810;
assign w8929 = ~w5812 & ~w8928;
assign w8930 = ~w5614 & ~w5616;
assign w8931 = ~w5617 & ~w8930;
assign w8932 = (w5598 & w5601) | (w5598 & w12880) | (w5601 & w12880);
assign w8933 = ~w5612 & ~w8932;
assign w8934 = ~w5540 & ~w5554;
assign w8935 = ~w5551 & ~w8934;
assign w8936 = ~w5573 & ~w5587;
assign w8937 = ~w5584 & ~w8936;
assign w8938 = ~w8935 & w8937;
assign w8939 = w8935 & ~w8937;
assign w8940 = ~w8938 & ~w8939;
assign w8941 = ~w8933 & ~w8940;
assign w8942 = ~w5612 & ~w8938;
assign w8943 = ~w8939 & w8942;
assign w8944 = ~w8932 & w8943;
assign w8945 = ~w8941 & ~w8944;
assign w8946 = (w5470 & w5506) | (w5470 & w12881) | (w5506 & w12881);
assign w8947 = ~w5513 & ~w8946;
assign w8948 = ~w5499 & ~w5503;
assign w8949 = ~w5496 & ~w8948;
assign w8950 = ~w5462 & ~w5465;
assign w8951 = ~w5468 & ~w8950;
assign w8952 = ~w8949 & w8951;
assign w8953 = w8949 & ~w8951;
assign w8954 = ~w8952 & ~w8953;
assign w8955 = ~w8947 & ~w8954;
assign w8956 = ~w5513 & ~w8952;
assign w8957 = ~w8953 & w8956;
assign w8958 = ~w8946 & w8957;
assign w8959 = ~w8955 & ~w8958;
assign w8960 = ~w8945 & w8959;
assign w8961 = w8945 & ~w8959;
assign w8962 = ~w8960 & ~w8961;
assign w8963 = ~w8931 & ~w8962;
assign w8964 = w8931 & w8962;
assign w8965 = ~w8963 & ~w8964;
assign w8966 = ~w5702 & ~w5795;
assign w8967 = ~w5796 & ~w8966;
assign w8968 = (w5653 & w5689) | (w5653 & w12882) | (w5689 & w12882);
assign w8969 = ~w5700 & ~w8968;
assign w8970 = ~w5682 & ~w5686;
assign w8971 = ~w5679 & ~w8970;
assign w8972 = ~w5645 & ~w5648;
assign w8973 = ~w5651 & ~w8972;
assign w8974 = ~w8971 & w8973;
assign w8975 = w8971 & ~w8973;
assign w8976 = ~w8974 & ~w8975;
assign w8977 = ~w8969 & ~w8976;
assign w8978 = ~w5700 & ~w8974;
assign w8979 = ~w8975 & w8978;
assign w8980 = ~w8968 & w8979;
assign w8981 = ~w8977 & ~w8980;
assign w8982 = (w5735 & w5771) | (w5735 & w12883) | (w5771 & w12883);
assign w8983 = ~w5778 & ~w8982;
assign w8984 = ~w5764 & ~w5768;
assign w8985 = ~w5761 & ~w8984;
assign w8986 = ~w5727 & ~w5730;
assign w8987 = ~w5733 & ~w8986;
assign w8988 = ~w8985 & w8987;
assign w8989 = w8985 & ~w8987;
assign w8990 = ~w8988 & ~w8989;
assign w8991 = ~w8983 & ~w8990;
assign w8992 = ~w5778 & ~w8988;
assign w8993 = ~w8989 & w8992;
assign w8994 = ~w8982 & w8993;
assign w8995 = ~w8991 & ~w8994;
assign w8996 = ~w8981 & w8995;
assign w8997 = w8981 & ~w8995;
assign w8998 = ~w8996 & ~w8997;
assign w8999 = ~w8967 & ~w8998;
assign w9000 = w8967 & w8998;
assign w9001 = ~w8999 & ~w9000;
assign w9002 = ~w8965 & w9001;
assign w9003 = w8965 & ~w9001;
assign w9004 = ~w9002 & ~w9003;
assign w9005 = ~w8929 & ~w9004;
assign w9006 = w8929 & w9004;
assign w9007 = ~w9005 & ~w9006;
assign w9008 = ~w8927 & w9007;
assign w9009 = w8927 & ~w9007;
assign w9010 = ~w9008 & ~w9009;
assign w9011 = ~w8847 & ~w9010;
assign w9012 = w8847 & w9010;
assign w9013 = ~w9011 & ~w9012;
assign w9014 = ~w8845 & w9013;
assign w9015 = w8845 & ~w9013;
assign w9016 = ~w9014 & ~w9015;
assign w9017 = ~w8677 & ~w9016;
assign w9018 = w8677 & w9016;
assign w9019 = ~w9017 & ~w9018;
assign w9020 = ~w7412 & ~w8199;
assign w9021 = ~w8201 & ~w9020;
assign w9022 = ~w7405 & ~w7408;
assign w9023 = ~w7409 & ~w9022;
assign w9024 = ~w7399 & ~w7402;
assign w9025 = ~w7403 & ~w9024;
assign w9026 = ~w7393 & ~w7395;
assign w9027 = ~w7396 & ~w9026;
assign w9028 = (w7377 & w7380) | (w7377 & w12884) | (w7380 & w12884);
assign w9029 = ~w7391 & ~w9028;
assign w9030 = ~w7243 & ~w7257;
assign w9031 = ~w7254 & ~w9030;
assign w9032 = ~w7276 & ~w7290;
assign w9033 = ~w7287 & ~w9032;
assign w9034 = ~w9031 & w9033;
assign w9035 = w9031 & ~w9033;
assign w9036 = ~w9034 & ~w9035;
assign w9037 = ~w9029 & ~w9036;
assign w9038 = ~w7391 & ~w9034;
assign w9039 = ~w9035 & w9038;
assign w9040 = ~w9028 & w9039;
assign w9041 = ~w9037 & ~w9040;
assign w9042 = (w7356 & w7359) | (w7356 & w12885) | (w7359 & w12885);
assign w9043 = ~w7366 & ~w9042;
assign w9044 = ~w7174 & ~w7188;
assign w9045 = ~w7185 & ~w9044;
assign w9046 = ~w7207 & ~w7221;
assign w9047 = ~w7218 & ~w9046;
assign w9048 = ~w9045 & w9047;
assign w9049 = w9045 & ~w9047;
assign w9050 = ~w9048 & ~w9049;
assign w9051 = ~w9043 & ~w9050;
assign w9052 = ~w7366 & ~w9048;
assign w9053 = ~w9049 & w9052;
assign w9054 = ~w9042 & w9053;
assign w9055 = ~w9051 & ~w9054;
assign w9056 = ~w9041 & w9055;
assign w9057 = w9041 & ~w9055;
assign w9058 = ~w9056 & ~w9057;
assign w9059 = ~w9027 & ~w9058;
assign w9060 = w9027 & w9058;
assign w9061 = ~w9059 & ~w9060;
assign w9062 = ~w7324 & ~w7343;
assign w9063 = ~w7344 & ~w9062;
assign w9064 = (w7308 & w7311) | (w7308 & w12886) | (w7311 & w12886);
assign w9065 = ~w7322 & ~w9064;
assign w9066 = ~w7102 & ~w7116;
assign w9067 = ~w7113 & ~w9066;
assign w9068 = ~w7135 & ~w7149;
assign w9069 = ~w7146 & ~w9068;
assign w9070 = ~w9067 & w9069;
assign w9071 = w9067 & ~w9069;
assign w9072 = ~w9070 & ~w9071;
assign w9073 = ~w9065 & ~w9072;
assign w9074 = ~w7322 & ~w9070;
assign w9075 = ~w9071 & w9074;
assign w9076 = ~w9064 & w9075;
assign w9077 = ~w9073 & ~w9076;
assign w9078 = (w7326 & w7329) | (w7326 & w12887) | (w7329 & w12887);
assign w9079 = ~w7336 & ~w9078;
assign w9080 = ~w7033 & ~w7047;
assign w9081 = ~w7044 & ~w9080;
assign w9082 = ~w7066 & ~w7080;
assign w9083 = ~w7077 & ~w9082;
assign w9084 = ~w9081 & w9083;
assign w9085 = w9081 & ~w9083;
assign w9086 = ~w9084 & ~w9085;
assign w9087 = ~w9079 & ~w9086;
assign w9088 = ~w7336 & ~w9084;
assign w9089 = ~w9085 & w9088;
assign w9090 = ~w9078 & w9089;
assign w9091 = ~w9087 & ~w9090;
assign w9092 = ~w9077 & w9091;
assign w9093 = w9077 & ~w9091;
assign w9094 = ~w9092 & ~w9093;
assign w9095 = ~w9063 & ~w9094;
assign w9096 = w9063 & w9094;
assign w9097 = ~w9095 & ~w9096;
assign w9098 = ~w9061 & w9097;
assign w9099 = w9061 & ~w9097;
assign w9100 = ~w9098 & ~w9099;
assign w9101 = ~w9025 & ~w9100;
assign w9102 = w9025 & w9100;
assign w9103 = ~w9101 & ~w9102;
assign w9104 = ~w6815 & ~w7005;
assign w9105 = ~w7007 & ~w9104;
assign w9106 = ~w6809 & ~w6811;
assign w9107 = ~w6812 & ~w9106;
assign w9108 = (w6793 & w6796) | (w6793 & w12888) | (w6796 & w12888);
assign w9109 = ~w6807 & ~w9108;
assign w9110 = ~w6735 & ~w6749;
assign w9111 = ~w6746 & ~w9110;
assign w9112 = ~w6768 & ~w6782;
assign w9113 = ~w6779 & ~w9112;
assign w9114 = ~w9111 & w9113;
assign w9115 = w9111 & ~w9113;
assign w9116 = ~w9114 & ~w9115;
assign w9117 = ~w9109 & ~w9116;
assign w9118 = ~w6807 & ~w9114;
assign w9119 = ~w9115 & w9118;
assign w9120 = ~w9108 & w9119;
assign w9121 = ~w9117 & ~w9120;
assign w9122 = (w6665 & w6701) | (w6665 & w12889) | (w6701 & w12889);
assign w9123 = ~w6708 & ~w9122;
assign w9124 = ~w6694 & ~w6698;
assign w9125 = ~w6691 & ~w9124;
assign w9126 = ~w6657 & ~w6660;
assign w9127 = ~w6663 & ~w9126;
assign w9128 = ~w9125 & w9127;
assign w9129 = w9125 & ~w9127;
assign w9130 = ~w9128 & ~w9129;
assign w9131 = ~w9123 & ~w9130;
assign w9132 = ~w6708 & ~w9128;
assign w9133 = ~w9129 & w9132;
assign w9134 = ~w9122 & w9133;
assign w9135 = ~w9131 & ~w9134;
assign w9136 = ~w9121 & w9135;
assign w9137 = w9121 & ~w9135;
assign w9138 = ~w9136 & ~w9137;
assign w9139 = ~w9107 & ~w9138;
assign w9140 = w9107 & w9138;
assign w9141 = ~w9139 & ~w9140;
assign w9142 = ~w6897 & ~w6990;
assign w9143 = ~w6991 & ~w9142;
assign w9144 = (w6848 & w6884) | (w6848 & w12890) | (w6884 & w12890);
assign w9145 = ~w6895 & ~w9144;
assign w9146 = ~w6877 & ~w6881;
assign w9147 = ~w6874 & ~w9146;
assign w9148 = ~w6840 & ~w6843;
assign w9149 = ~w6846 & ~w9148;
assign w9150 = ~w9147 & w9149;
assign w9151 = w9147 & ~w9149;
assign w9152 = ~w9150 & ~w9151;
assign w9153 = ~w9145 & ~w9152;
assign w9154 = ~w6895 & ~w9150;
assign w9155 = ~w9151 & w9154;
assign w9156 = ~w9144 & w9155;
assign w9157 = ~w9153 & ~w9156;
assign w9158 = (w6930 & w6966) | (w6930 & w12891) | (w6966 & w12891);
assign w9159 = ~w6973 & ~w9158;
assign w9160 = ~w6959 & ~w6963;
assign w9161 = ~w6956 & ~w9160;
assign w9162 = ~w6922 & ~w6925;
assign w9163 = ~w6928 & ~w9162;
assign w9164 = ~w9161 & w9163;
assign w9165 = w9161 & ~w9163;
assign w9166 = ~w9164 & ~w9165;
assign w9167 = ~w9159 & ~w9166;
assign w9168 = ~w6973 & ~w9164;
assign w9169 = ~w9165 & w9168;
assign w9170 = ~w9158 & w9169;
assign w9171 = ~w9167 & ~w9170;
assign w9172 = ~w9157 & w9171;
assign w9173 = w9157 & ~w9171;
assign w9174 = ~w9172 & ~w9173;
assign w9175 = ~w9143 & ~w9174;
assign w9176 = w9143 & w9174;
assign w9177 = ~w9175 & ~w9176;
assign w9178 = ~w9141 & w9177;
assign w9179 = w9141 & ~w9177;
assign w9180 = ~w9178 & ~w9179;
assign w9181 = ~w9105 & ~w9180;
assign w9182 = w9105 & w9180;
assign w9183 = ~w9181 & ~w9182;
assign w9184 = ~w9103 & w9183;
assign w9185 = w9103 & ~w9183;
assign w9186 = ~w9184 & ~w9185;
assign w9187 = ~w9023 & ~w9186;
assign w9188 = w9023 & w9186;
assign w9189 = ~w9187 & ~w9188;
assign w9190 = ~w7793 & ~w8182;
assign w9191 = ~w8183 & ~w9190;
assign w9192 = ~w7787 & ~w7790;
assign w9193 = ~w7791 & ~w9192;
assign w9194 = ~w7781 & ~w7783;
assign w9195 = ~w7784 & ~w9194;
assign w9196 = (w7765 & w7768) | (w7765 & w12892) | (w7768 & w12892);
assign w9197 = ~w7779 & ~w9196;
assign w9198 = ~w7682 & ~w7696;
assign w9199 = ~w7693 & ~w9198;
assign w9200 = ~w7715 & ~w7729;
assign w9201 = ~w7726 & ~w9200;
assign w9202 = ~w9199 & w9201;
assign w9203 = w9199 & ~w9201;
assign w9204 = ~w9202 & ~w9203;
assign w9205 = ~w9197 & ~w9204;
assign w9206 = ~w7779 & ~w9202;
assign w9207 = ~w9203 & w9206;
assign w9208 = ~w9196 & w9207;
assign w9209 = ~w9205 & ~w9208;
assign w9210 = (w7744 & w7747) | (w7744 & w12893) | (w7747 & w12893);
assign w9211 = ~w7754 & ~w9210;
assign w9212 = ~w7613 & ~w7627;
assign w9213 = ~w7624 & ~w9212;
assign w9214 = ~w7646 & ~w7660;
assign w9215 = ~w7657 & ~w9214;
assign w9216 = ~w9213 & w9215;
assign w9217 = w9213 & ~w9215;
assign w9218 = ~w9216 & ~w9217;
assign w9219 = ~w9211 & ~w9218;
assign w9220 = ~w7754 & ~w9216;
assign w9221 = ~w9217 & w9220;
assign w9222 = ~w9210 & w9221;
assign w9223 = ~w9219 & ~w9222;
assign w9224 = ~w9209 & w9223;
assign w9225 = w9209 & ~w9223;
assign w9226 = ~w9224 & ~w9225;
assign w9227 = ~w9195 & ~w9226;
assign w9228 = w9195 & w9226;
assign w9229 = ~w9227 & ~w9228;
assign w9230 = ~w7494 & ~w7587;
assign w9231 = ~w7588 & ~w9230;
assign w9232 = (w7445 & w7481) | (w7445 & w12894) | (w7481 & w12894);
assign w9233 = ~w7492 & ~w9232;
assign w9234 = ~w7474 & ~w7478;
assign w9235 = ~w7471 & ~w9234;
assign w9236 = ~w7437 & ~w7440;
assign w9237 = ~w7443 & ~w9236;
assign w9238 = ~w9235 & w9237;
assign w9239 = w9235 & ~w9237;
assign w9240 = ~w9238 & ~w9239;
assign w9241 = ~w9233 & ~w9240;
assign w9242 = ~w7492 & ~w9238;
assign w9243 = ~w9239 & w9242;
assign w9244 = ~w9232 & w9243;
assign w9245 = ~w9241 & ~w9244;
assign w9246 = (w7527 & w7563) | (w7527 & w12895) | (w7563 & w12895);
assign w9247 = ~w7570 & ~w9246;
assign w9248 = ~w7556 & ~w7560;
assign w9249 = ~w7553 & ~w9248;
assign w9250 = ~w7519 & ~w7522;
assign w9251 = ~w7525 & ~w9250;
assign w9252 = ~w9249 & w9251;
assign w9253 = w9249 & ~w9251;
assign w9254 = ~w9252 & ~w9253;
assign w9255 = ~w9247 & ~w9254;
assign w9256 = ~w7570 & ~w9252;
assign w9257 = ~w9253 & w9256;
assign w9258 = ~w9246 & w9257;
assign w9259 = ~w9255 & ~w9258;
assign w9260 = ~w9245 & w9259;
assign w9261 = w9245 & ~w9259;
assign w9262 = ~w9260 & ~w9261;
assign w9263 = ~w9231 & ~w9262;
assign w9264 = w9231 & w9262;
assign w9265 = ~w9263 & ~w9264;
assign w9266 = ~w9229 & w9265;
assign w9267 = w9229 & ~w9265;
assign w9268 = ~w9266 & ~w9267;
assign w9269 = ~w9193 & ~w9268;
assign w9270 = w9193 & w9268;
assign w9271 = ~w9269 & ~w9270;
assign w9272 = ~w7975 & ~w8165;
assign w9273 = ~w8167 & ~w9272;
assign w9274 = ~w7970 & ~w7972;
assign w9275 = ~w7973 & ~w9274;
assign w9276 = (w7954 & w7957) | (w7954 & w12896) | (w7957 & w12896);
assign w9277 = ~w7968 & ~w9276;
assign w9278 = ~w7896 & ~w7910;
assign w9279 = ~w7907 & ~w9278;
assign w9280 = ~w7929 & ~w7943;
assign w9281 = ~w7940 & ~w9280;
assign w9282 = ~w9279 & w9281;
assign w9283 = w9279 & ~w9281;
assign w9284 = ~w9282 & ~w9283;
assign w9285 = ~w9277 & ~w9284;
assign w9286 = ~w7968 & ~w9282;
assign w9287 = ~w9283 & w9286;
assign w9288 = ~w9276 & w9287;
assign w9289 = ~w9285 & ~w9288;
assign w9290 = (w7826 & w7862) | (w7826 & w12897) | (w7862 & w12897);
assign w9291 = ~w7869 & ~w9290;
assign w9292 = ~w7855 & ~w7859;
assign w9293 = ~w7852 & ~w9292;
assign w9294 = ~w7818 & ~w7821;
assign w9295 = ~w7824 & ~w9294;
assign w9296 = ~w9293 & w9295;
assign w9297 = w9293 & ~w9295;
assign w9298 = ~w9296 & ~w9297;
assign w9299 = ~w9291 & ~w9298;
assign w9300 = ~w7869 & ~w9296;
assign w9301 = ~w9297 & w9300;
assign w9302 = ~w9290 & w9301;
assign w9303 = ~w9299 & ~w9302;
assign w9304 = ~w9289 & w9303;
assign w9305 = w9289 & ~w9303;
assign w9306 = ~w9304 & ~w9305;
assign w9307 = ~w9275 & ~w9306;
assign w9308 = w9275 & w9306;
assign w9309 = ~w9307 & ~w9308;
assign w9310 = ~w8057 & ~w8150;
assign w9311 = ~w8151 & ~w9310;
assign w9312 = (w8008 & w8044) | (w8008 & w12898) | (w8044 & w12898);
assign w9313 = ~w8055 & ~w9312;
assign w9314 = ~w8037 & ~w8041;
assign w9315 = ~w8034 & ~w9314;
assign w9316 = ~w8000 & ~w8003;
assign w9317 = ~w8006 & ~w9316;
assign w9318 = ~w9315 & w9317;
assign w9319 = w9315 & ~w9317;
assign w9320 = ~w9318 & ~w9319;
assign w9321 = ~w9313 & ~w9320;
assign w9322 = ~w8055 & ~w9318;
assign w9323 = ~w9319 & w9322;
assign w9324 = ~w9312 & w9323;
assign w9325 = ~w9321 & ~w9324;
assign w9326 = (w8090 & w8126) | (w8090 & w12899) | (w8126 & w12899);
assign w9327 = ~w8133 & ~w9326;
assign w9328 = ~w8119 & ~w8123;
assign w9329 = ~w8116 & ~w9328;
assign w9330 = ~w8082 & ~w8085;
assign w9331 = ~w8088 & ~w9330;
assign w9332 = ~w9329 & w9331;
assign w9333 = w9329 & ~w9331;
assign w9334 = ~w9332 & ~w9333;
assign w9335 = ~w9327 & ~w9334;
assign w9336 = ~w8133 & ~w9332;
assign w9337 = ~w9333 & w9336;
assign w9338 = ~w9326 & w9337;
assign w9339 = ~w9335 & ~w9338;
assign w9340 = ~w9325 & w9339;
assign w9341 = w9325 & ~w9339;
assign w9342 = ~w9340 & ~w9341;
assign w9343 = ~w9311 & ~w9342;
assign w9344 = w9311 & w9342;
assign w9345 = ~w9343 & ~w9344;
assign w9346 = ~w9309 & w9345;
assign w9347 = w9309 & ~w9345;
assign w9348 = ~w9346 & ~w9347;
assign w9349 = ~w9273 & ~w9348;
assign w9350 = w9273 & w9348;
assign w9351 = ~w9349 & ~w9350;
assign w9352 = ~w9271 & w9351;
assign w9353 = w9271 & ~w9351;
assign w9354 = ~w9352 & ~w9353;
assign w9355 = ~w9191 & ~w9354;
assign w9356 = w9191 & w9354;
assign w9357 = ~w9355 & ~w9356;
assign w9358 = ~w9189 & w9357;
assign w9359 = w9189 & ~w9357;
assign w9360 = ~w9358 & ~w9359;
assign w9361 = ~w9021 & ~w9360;
assign w9362 = w9021 & w9360;
assign w9363 = ~w9361 & ~w9362;
assign w9364 = ~w9019 & w9363;
assign w9365 = w9019 & ~w9363;
assign w9366 = ~w9364 & ~w9365;
assign w9367 = ~w8675 & ~w9366;
assign w9368 = w8675 & w9366;
assign w9369 = ~w9367 & ~w9368;
assign w9370 = ~w8673 & w9369;
assign w9371 = w8673 & ~w9369;
assign w9372 = ~w9370 & ~w9371;
assign w9373 = ~w8256 & ~w9372;
assign w9374 = w8256 & w9372;
assign w9375 = ~w9373 & ~w9374;
assign w9376 = ~w3155 & ~w3158;
assign w9377 = ~w3159 & ~w9376;
assign w9378 = ~w3149 & ~w3152;
assign w9379 = ~w3153 & ~w9378;
assign w9380 = ~w3142 & ~w3145;
assign w9381 = ~w3146 & ~w9380;
assign w9382 = ~w3136 & ~w3139;
assign w9383 = ~w3140 & ~w9382;
assign w9384 = ~w3131 & ~w3133;
assign w9385 = ~w3134 & ~w9384;
assign w9386 = (w3115 & w3118) | (w3115 & w13550) | (w3118 & w13550);
assign w9387 = ~w3129 & ~w9386;
assign w9388 = ~w1588 & ~w1602;
assign w9389 = ~w1599 & ~w9388;
assign w9390 = ~w1621 & ~w1632;
assign w9391 = ~w1635 & ~w9390;
assign w9392 = ~w9389 & w9391;
assign w9393 = w9389 & ~w9391;
assign w9394 = ~w9392 & ~w9393;
assign w9395 = ~w9387 & ~w9394;
assign w9396 = ~w3129 & ~w9392;
assign w9397 = ~w9393 & w9396;
assign w9398 = ~w9386 & w9397;
assign w9399 = ~w9395 & ~w9398;
assign w9400 = (w3094 & w3097) | (w3094 & w13551) | (w3097 & w13551);
assign w9401 = ~w3104 & ~w9400;
assign w9402 = ~w1657 & ~w1671;
assign w9403 = ~w1668 & ~w9402;
assign w9404 = ~w1690 & ~w1704;
assign w9405 = ~w1701 & ~w9404;
assign w9406 = ~w9403 & w9405;
assign w9407 = w9403 & ~w9405;
assign w9408 = ~w9406 & ~w9407;
assign w9409 = ~w9401 & ~w9408;
assign w9410 = ~w3104 & ~w9406;
assign w9411 = ~w9407 & w9410;
assign w9412 = ~w9400 & w9411;
assign w9413 = ~w9409 & ~w9412;
assign w9414 = ~w9399 & w9413;
assign w9415 = w9399 & ~w9413;
assign w9416 = ~w9414 & ~w9415;
assign w9417 = ~w9385 & ~w9416;
assign w9418 = w9385 & w9416;
assign w9419 = ~w9417 & ~w9418;
assign w9420 = ~w3062 & ~w3081;
assign w9421 = ~w3082 & ~w9420;
assign w9422 = (w3046 & w3049) | (w3046 & w13552) | (w3049 & w13552);
assign w9423 = ~w3060 & ~w9422;
assign w9424 = ~w1798 & ~w1812;
assign w9425 = ~w1809 & ~w9424;
assign w9426 = ~w1831 & ~w1845;
assign w9427 = ~w1842 & ~w9426;
assign w9428 = ~w9425 & w9427;
assign w9429 = w9425 & ~w9427;
assign w9430 = ~w9428 & ~w9429;
assign w9431 = ~w9423 & ~w9430;
assign w9432 = ~w3060 & ~w9428;
assign w9433 = ~w9429 & w9432;
assign w9434 = ~w9422 & w9433;
assign w9435 = ~w9431 & ~w9434;
assign w9436 = (w3064 & w3067) | (w3064 & w13553) | (w3067 & w13553);
assign w9437 = ~w3074 & ~w9436;
assign w9438 = ~w1729 & ~w1743;
assign w9439 = ~w1740 & ~w9438;
assign w9440 = ~w1762 & ~w1776;
assign w9441 = ~w1773 & ~w9440;
assign w9442 = ~w9439 & w9441;
assign w9443 = w9439 & ~w9441;
assign w9444 = ~w9442 & ~w9443;
assign w9445 = ~w9437 & ~w9444;
assign w9446 = ~w3074 & ~w9442;
assign w9447 = ~w9443 & w9446;
assign w9448 = ~w9436 & w9447;
assign w9449 = ~w9445 & ~w9448;
assign w9450 = ~w9435 & w9449;
assign w9451 = w9435 & ~w9449;
assign w9452 = ~w9450 & ~w9451;
assign w9453 = ~w9421 & ~w9452;
assign w9454 = w9421 & w9452;
assign w9455 = ~w9453 & ~w9454;
assign w9456 = ~w9419 & w9455;
assign w9457 = w9419 & ~w9455;
assign w9458 = ~w9456 & ~w9457;
assign w9459 = ~w9383 & ~w9458;
assign w9460 = w9383 & w9458;
assign w9461 = ~w9459 & ~w9460;
assign w9462 = ~w2985 & ~w3031;
assign w9463 = ~w3033 & ~w9462;
assign w9464 = ~w2980 & ~w2982;
assign w9465 = ~w2983 & ~w9464;
assign w9466 = (w2964 & w2967) | (w2964 & w13554) | (w2967 & w13554);
assign w9467 = ~w2978 & ~w9466;
assign w9468 = ~w2083 & ~w2097;
assign w9469 = ~w2094 & ~w9468;
assign w9470 = ~w2116 & ~w2130;
assign w9471 = ~w2127 & ~w9470;
assign w9472 = ~w9469 & w9471;
assign w9473 = w9469 & ~w9471;
assign w9474 = ~w9472 & ~w9473;
assign w9475 = ~w9467 & ~w9474;
assign w9476 = ~w2978 & ~w9472;
assign w9477 = ~w9473 & w9476;
assign w9478 = ~w9466 & w9477;
assign w9479 = ~w9475 & ~w9478;
assign w9480 = (w2943 & w2946) | (w2943 & w13555) | (w2946 & w13555);
assign w9481 = ~w2953 & ~w9480;
assign w9482 = ~w2014 & ~w2028;
assign w9483 = ~w2025 & ~w9482;
assign w9484 = ~w2047 & ~w2061;
assign w9485 = ~w2058 & ~w9484;
assign w9486 = ~w9483 & w9485;
assign w9487 = w9483 & ~w9485;
assign w9488 = ~w9486 & ~w9487;
assign w9489 = ~w9481 & ~w9488;
assign w9490 = ~w2953 & ~w9486;
assign w9491 = ~w9487 & w9490;
assign w9492 = ~w9480 & w9491;
assign w9493 = ~w9489 & ~w9492;
assign w9494 = ~w9479 & w9493;
assign w9495 = w9479 & ~w9493;
assign w9496 = ~w9494 & ~w9495;
assign w9497 = ~w9465 & ~w9496;
assign w9498 = w9465 & w9496;
assign w9499 = ~w9497 & ~w9498;
assign w9500 = ~w3003 & ~w3022;
assign w9501 = ~w3023 & ~w9500;
assign w9502 = (w2987 & w2990) | (w2987 & w13556) | (w2990 & w13556);
assign w9503 = ~w3001 & ~w9502;
assign w9504 = ~w1942 & ~w1956;
assign w9505 = ~w1953 & ~w9504;
assign w9506 = ~w1975 & ~w1989;
assign w9507 = ~w1986 & ~w9506;
assign w9508 = ~w9505 & w9507;
assign w9509 = w9505 & ~w9507;
assign w9510 = ~w9508 & ~w9509;
assign w9511 = ~w9503 & ~w9510;
assign w9512 = ~w3001 & ~w9508;
assign w9513 = ~w9509 & w9512;
assign w9514 = ~w9502 & w9513;
assign w9515 = ~w9511 & ~w9514;
assign w9516 = (w3005 & w3008) | (w3005 & w13557) | (w3008 & w13557);
assign w9517 = ~w3015 & ~w9516;
assign w9518 = ~w1873 & ~w1887;
assign w9519 = ~w1884 & ~w9518;
assign w9520 = ~w1906 & ~w1920;
assign w9521 = ~w1917 & ~w9520;
assign w9522 = ~w9519 & w9521;
assign w9523 = w9519 & ~w9521;
assign w9524 = ~w9522 & ~w9523;
assign w9525 = ~w9517 & ~w9524;
assign w9526 = ~w3015 & ~w9522;
assign w9527 = ~w9523 & w9526;
assign w9528 = ~w9516 & w9527;
assign w9529 = ~w9525 & ~w9528;
assign w9530 = ~w9515 & w9529;
assign w9531 = w9515 & ~w9529;
assign w9532 = ~w9530 & ~w9531;
assign w9533 = ~w9501 & ~w9532;
assign w9534 = w9501 & w9532;
assign w9535 = ~w9533 & ~w9534;
assign w9536 = ~w9499 & w9535;
assign w9537 = w9499 & ~w9535;
assign w9538 = ~w9536 & ~w9537;
assign w9539 = ~w9463 & ~w9538;
assign w9540 = w9463 & w9538;
assign w9541 = ~w9539 & ~w9540;
assign w9542 = ~w9461 & w9541;
assign w9543 = w9461 & ~w9541;
assign w9544 = ~w9542 & ~w9543;
assign w9545 = ~w9381 & ~w9544;
assign w9546 = w9381 & w9544;
assign w9547 = ~w9545 & ~w9546;
assign w9548 = ~w2826 & ~w2927;
assign w9549 = ~w2929 & ~w9548;
assign w9550 = ~w2820 & ~w2823;
assign w9551 = ~w2824 & ~w9550;
assign w9552 = ~w2815 & ~w2817;
assign w9553 = ~w2818 & ~w9552;
assign w9554 = (w2799 & w2802) | (w2799 & w13558) | (w2802 & w13558);
assign w9555 = ~w2813 & ~w9554;
assign w9556 = ~w2656 & ~w2670;
assign w9557 = ~w2667 & ~w9556;
assign w9558 = ~w2689 & ~w2703;
assign w9559 = ~w2700 & ~w9558;
assign w9560 = ~w9557 & w9559;
assign w9561 = w9557 & ~w9559;
assign w9562 = ~w9560 & ~w9561;
assign w9563 = ~w9555 & ~w9562;
assign w9564 = ~w2813 & ~w9560;
assign w9565 = ~w9561 & w9564;
assign w9566 = ~w9554 & w9565;
assign w9567 = ~w9563 & ~w9566;
assign w9568 = (w2778 & w2781) | (w2778 & w13559) | (w2781 & w13559);
assign w9569 = ~w2788 & ~w9568;
assign w9570 = ~w2587 & ~w2601;
assign w9571 = ~w2598 & ~w9570;
assign w9572 = ~w2620 & ~w2634;
assign w9573 = ~w2631 & ~w9572;
assign w9574 = ~w9571 & w9573;
assign w9575 = w9571 & ~w9573;
assign w9576 = ~w9574 & ~w9575;
assign w9577 = ~w9569 & ~w9576;
assign w9578 = ~w2788 & ~w9574;
assign w9579 = ~w9575 & w9578;
assign w9580 = ~w9568 & w9579;
assign w9581 = ~w9577 & ~w9580;
assign w9582 = ~w9567 & w9581;
assign w9583 = w9567 & ~w9581;
assign w9584 = ~w9582 & ~w9583;
assign w9585 = ~w9553 & ~w9584;
assign w9586 = w9553 & w9584;
assign w9587 = ~w9585 & ~w9586;
assign w9588 = ~w2746 & ~w2765;
assign w9589 = ~w2766 & ~w9588;
assign w9590 = (w2730 & w2733) | (w2730 & w13560) | (w2733 & w13560);
assign w9591 = ~w2744 & ~w9590;
assign w9592 = ~w2515 & ~w2529;
assign w9593 = ~w2526 & ~w9592;
assign w9594 = ~w2548 & ~w2562;
assign w9595 = ~w2559 & ~w9594;
assign w9596 = ~w9593 & w9595;
assign w9597 = w9593 & ~w9595;
assign w9598 = ~w9596 & ~w9597;
assign w9599 = ~w9591 & ~w9598;
assign w9600 = ~w2744 & ~w9596;
assign w9601 = ~w9597 & w9600;
assign w9602 = ~w9590 & w9601;
assign w9603 = ~w9599 & ~w9602;
assign w9604 = (w2748 & w2751) | (w2748 & w13561) | (w2751 & w13561);
assign w9605 = ~w2758 & ~w9604;
assign w9606 = ~w2446 & ~w2460;
assign w9607 = ~w2457 & ~w9606;
assign w9608 = ~w2479 & ~w2493;
assign w9609 = ~w2490 & ~w9608;
assign w9610 = ~w9607 & w9609;
assign w9611 = w9607 & ~w9609;
assign w9612 = ~w9610 & ~w9611;
assign w9613 = ~w9605 & ~w9612;
assign w9614 = ~w2758 & ~w9610;
assign w9615 = ~w9611 & w9614;
assign w9616 = ~w9604 & w9615;
assign w9617 = ~w9613 & ~w9616;
assign w9618 = ~w9603 & w9617;
assign w9619 = w9603 & ~w9617;
assign w9620 = ~w9618 & ~w9619;
assign w9621 = ~w9589 & ~w9620;
assign w9622 = w9589 & w9620;
assign w9623 = ~w9621 & ~w9622;
assign w9624 = ~w9587 & w9623;
assign w9625 = w9587 & ~w9623;
assign w9626 = ~w9624 & ~w9625;
assign w9627 = ~w9551 & ~w9626;
assign w9628 = w9551 & w9626;
assign w9629 = ~w9627 & ~w9628;
assign w9630 = ~w2870 & ~w2916;
assign w9631 = ~w2918 & ~w9630;
assign w9632 = ~w2865 & ~w2867;
assign w9633 = ~w2868 & ~w9632;
assign w9634 = (w2849 & w2852) | (w2849 & w13562) | (w2852 & w13562);
assign w9635 = ~w2863 & ~w9634;
assign w9636 = ~w2371 & ~w2385;
assign w9637 = ~w2382 & ~w9636;
assign w9638 = ~w2404 & ~w2418;
assign w9639 = ~w2415 & ~w9638;
assign w9640 = ~w9637 & w9639;
assign w9641 = w9637 & ~w9639;
assign w9642 = ~w9640 & ~w9641;
assign w9643 = ~w9635 & ~w9642;
assign w9644 = ~w2863 & ~w9640;
assign w9645 = ~w9641 & w9644;
assign w9646 = ~w9634 & w9645;
assign w9647 = ~w9643 & ~w9646;
assign w9648 = (w2828 & w2831) | (w2828 & w13563) | (w2831 & w13563);
assign w9649 = ~w2838 & ~w9648;
assign w9650 = ~w2302 & ~w2316;
assign w9651 = ~w2313 & ~w9650;
assign w9652 = ~w2335 & ~w2349;
assign w9653 = ~w2346 & ~w9652;
assign w9654 = ~w9651 & w9653;
assign w9655 = w9651 & ~w9653;
assign w9656 = ~w9654 & ~w9655;
assign w9657 = ~w9649 & ~w9656;
assign w9658 = ~w2838 & ~w9654;
assign w9659 = ~w9655 & w9658;
assign w9660 = ~w9648 & w9659;
assign w9661 = ~w9657 & ~w9660;
assign w9662 = ~w9647 & w9661;
assign w9663 = w9647 & ~w9661;
assign w9664 = ~w9662 & ~w9663;
assign w9665 = ~w9633 & ~w9664;
assign w9666 = w9633 & w9664;
assign w9667 = ~w9665 & ~w9666;
assign w9668 = ~w2888 & ~w2907;
assign w9669 = ~w2908 & ~w9668;
assign w9670 = (w2872 & w2875) | (w2872 & w13564) | (w2875 & w13564);
assign w9671 = ~w2886 & ~w9670;
assign w9672 = ~w2230 & ~w2244;
assign w9673 = ~w2241 & ~w9672;
assign w9674 = ~w2263 & ~w2277;
assign w9675 = ~w2274 & ~w9674;
assign w9676 = ~w9673 & w9675;
assign w9677 = w9673 & ~w9675;
assign w9678 = ~w9676 & ~w9677;
assign w9679 = ~w9671 & ~w9678;
assign w9680 = ~w2886 & ~w9676;
assign w9681 = ~w9677 & w9680;
assign w9682 = ~w9670 & w9681;
assign w9683 = ~w9679 & ~w9682;
assign w9684 = (w2890 & w2893) | (w2890 & w13565) | (w2893 & w13565);
assign w9685 = ~w2900 & ~w9684;
assign w9686 = ~w2161 & ~w2175;
assign w9687 = ~w2172 & ~w9686;
assign w9688 = ~w2194 & ~w2208;
assign w9689 = ~w2205 & ~w9688;
assign w9690 = ~w9687 & w9689;
assign w9691 = w9687 & ~w9689;
assign w9692 = ~w9690 & ~w9691;
assign w9693 = ~w9685 & ~w9692;
assign w9694 = ~w2900 & ~w9690;
assign w9695 = ~w9691 & w9694;
assign w9696 = ~w9684 & w9695;
assign w9697 = ~w9693 & ~w9696;
assign w9698 = ~w9683 & w9697;
assign w9699 = w9683 & ~w9697;
assign w9700 = ~w9698 & ~w9699;
assign w9701 = ~w9669 & ~w9700;
assign w9702 = w9669 & w9700;
assign w9703 = ~w9701 & ~w9702;
assign w9704 = ~w9667 & w9703;
assign w9705 = w9667 & ~w9703;
assign w9706 = ~w9704 & ~w9705;
assign w9707 = ~w9631 & ~w9706;
assign w9708 = w9631 & w9706;
assign w9709 = ~w9707 & ~w9708;
assign w9710 = ~w9629 & w9709;
assign w9711 = w9629 & ~w9709;
assign w9712 = ~w9710 & ~w9711;
assign w9713 = ~w9549 & ~w9712;
assign w9714 = w9549 & w9712;
assign w9715 = ~w9713 & ~w9714;
assign w9716 = ~w9547 & w9715;
assign w9717 = w9547 & ~w9715;
assign w9718 = ~w9716 & ~w9717;
assign w9719 = ~w9379 & ~w9718;
assign w9720 = w9379 & w9718;
assign w9721 = ~w9719 & ~w9720;
assign w9722 = ~w777 & ~w1563;
assign w9723 = ~w1565 & ~w9722;
assign w9724 = ~w770 & ~w773;
assign w9725 = ~w774 & ~w9724;
assign w9726 = ~w764 & ~w767;
assign w9727 = ~w768 & ~w9726;
assign w9728 = ~w759 & ~w761;
assign w9729 = ~w762 & ~w9728;
assign w9730 = (w743 & w746) | (w743 & w13566) | (w746 & w13566);
assign w9731 = ~w757 & ~w9730;
assign w9732 = ~w608 & ~w622;
assign w9733 = ~w619 & ~w9732;
assign w9734 = ~w641 & ~w655;
assign w9735 = ~w652 & ~w9734;
assign w9736 = ~w9733 & w9735;
assign w9737 = w9733 & ~w9735;
assign w9738 = ~w9736 & ~w9737;
assign w9739 = ~w9731 & ~w9738;
assign w9740 = ~w757 & ~w9736;
assign w9741 = ~w9737 & w9740;
assign w9742 = ~w9730 & w9741;
assign w9743 = ~w9739 & ~w9742;
assign w9744 = (w722 & w725) | (w722 & w13567) | (w725 & w13567);
assign w9745 = ~w732 & ~w9744;
assign w9746 = ~w539 & ~w553;
assign w9747 = ~w550 & ~w9746;
assign w9748 = ~w572 & ~w586;
assign w9749 = ~w583 & ~w9748;
assign w9750 = ~w9747 & w9749;
assign w9751 = w9747 & ~w9749;
assign w9752 = ~w9750 & ~w9751;
assign w9753 = ~w9745 & ~w9752;
assign w9754 = ~w732 & ~w9750;
assign w9755 = ~w9751 & w9754;
assign w9756 = ~w9744 & w9755;
assign w9757 = ~w9753 & ~w9756;
assign w9758 = ~w9743 & w9757;
assign w9759 = w9743 & ~w9757;
assign w9760 = ~w9758 & ~w9759;
assign w9761 = ~w9729 & ~w9760;
assign w9762 = w9729 & w9760;
assign w9763 = ~w9761 & ~w9762;
assign w9764 = ~w690 & ~w709;
assign w9765 = ~w710 & ~w9764;
assign w9766 = (w674 & w677) | (w674 & w13568) | (w677 & w13568);
assign w9767 = ~w688 & ~w9766;
assign w9768 = ~w467 & ~w481;
assign w9769 = ~w478 & ~w9768;
assign w9770 = ~w500 & ~w514;
assign w9771 = ~w511 & ~w9770;
assign w9772 = ~w9769 & w9771;
assign w9773 = w9769 & ~w9771;
assign w9774 = ~w9772 & ~w9773;
assign w9775 = ~w9767 & ~w9774;
assign w9776 = ~w688 & ~w9772;
assign w9777 = ~w9773 & w9776;
assign w9778 = ~w9766 & w9777;
assign w9779 = ~w9775 & ~w9778;
assign w9780 = (w692 & w695) | (w692 & w13569) | (w695 & w13569);
assign w9781 = ~w702 & ~w9780;
assign w9782 = ~w398 & ~w412;
assign w9783 = ~w409 & ~w9782;
assign w9784 = ~w431 & ~w445;
assign w9785 = ~w442 & ~w9784;
assign w9786 = ~w9783 & w9785;
assign w9787 = w9783 & ~w9785;
assign w9788 = ~w9786 & ~w9787;
assign w9789 = ~w9781 & ~w9788;
assign w9790 = ~w702 & ~w9786;
assign w9791 = ~w9787 & w9790;
assign w9792 = ~w9780 & w9791;
assign w9793 = ~w9789 & ~w9792;
assign w9794 = ~w9779 & w9793;
assign w9795 = w9779 & ~w9793;
assign w9796 = ~w9794 & ~w9795;
assign w9797 = ~w9765 & ~w9796;
assign w9798 = w9765 & w9796;
assign w9799 = ~w9797 & ~w9798;
assign w9800 = ~w9763 & w9799;
assign w9801 = w9763 & ~w9799;
assign w9802 = ~w9800 & ~w9801;
assign w9803 = ~w9727 & ~w9802;
assign w9804 = w9727 & w9802;
assign w9805 = ~w9803 & ~w9804;
assign w9806 = ~w181 & ~w371;
assign w9807 = ~w373 & ~w9806;
assign w9808 = ~w176 & ~w178;
assign w9809 = ~w179 & ~w9808;
assign w9810 = (w160 & w163) | (w160 & w13570) | (w163 & w13570);
assign w9811 = ~w174 & ~w9810;
assign w9812 = ~w102 & ~w116;
assign w9813 = ~w113 & ~w9812;
assign w9814 = ~w135 & ~w149;
assign w9815 = ~w146 & ~w9814;
assign w9816 = ~w9813 & w9815;
assign w9817 = w9813 & ~w9815;
assign w9818 = ~w9816 & ~w9817;
assign w9819 = ~w9811 & ~w9818;
assign w9820 = ~w174 & ~w9816;
assign w9821 = ~w9817 & w9820;
assign w9822 = ~w9810 & w9821;
assign w9823 = ~w9819 & ~w9822;
assign w9824 = (w32 & w68) | (w32 & w13571) | (w68 & w13571);
assign w9825 = ~w75 & ~w9824;
assign w9826 = ~w61 & ~w65;
assign w9827 = ~w58 & ~w9826;
assign w9828 = ~w24 & ~w27;
assign w9829 = ~w30 & ~w9828;
assign w9830 = ~w9827 & w9829;
assign w9831 = w9827 & ~w9829;
assign w9832 = ~w9830 & ~w9831;
assign w9833 = ~w9825 & ~w9832;
assign w9834 = ~w75 & ~w9830;
assign w9835 = ~w9831 & w9834;
assign w9836 = ~w9824 & w9835;
assign w9837 = ~w9833 & ~w9836;
assign w9838 = ~w9823 & w9837;
assign w9839 = w9823 & ~w9837;
assign w9840 = ~w9838 & ~w9839;
assign w9841 = ~w9809 & ~w9840;
assign w9842 = w9809 & w9840;
assign w9843 = ~w9841 & ~w9842;
assign w9844 = ~w263 & ~w356;
assign w9845 = ~w357 & ~w9844;
assign w9846 = (w214 & w250) | (w214 & w13572) | (w250 & w13572);
assign w9847 = ~w261 & ~w9846;
assign w9848 = ~w243 & ~w247;
assign w9849 = ~w240 & ~w9848;
assign w9850 = ~w206 & ~w209;
assign w9851 = ~w212 & ~w9850;
assign w9852 = ~w9849 & w9851;
assign w9853 = w9849 & ~w9851;
assign w9854 = ~w9852 & ~w9853;
assign w9855 = ~w9847 & ~w9854;
assign w9856 = ~w261 & ~w9852;
assign w9857 = ~w9853 & w9856;
assign w9858 = ~w9846 & w9857;
assign w9859 = ~w9855 & ~w9858;
assign w9860 = (w296 & w332) | (w296 & w13573) | (w332 & w13573);
assign w9861 = ~w339 & ~w9860;
assign w9862 = ~w325 & ~w329;
assign w9863 = ~w322 & ~w9862;
assign w9864 = ~w288 & ~w291;
assign w9865 = ~w294 & ~w9864;
assign w9866 = ~w9863 & w9865;
assign w9867 = w9863 & ~w9865;
assign w9868 = ~w9866 & ~w9867;
assign w9869 = ~w9861 & ~w9868;
assign w9870 = ~w339 & ~w9866;
assign w9871 = ~w9867 & w9870;
assign w9872 = ~w9860 & w9871;
assign w9873 = ~w9869 & ~w9872;
assign w9874 = ~w9859 & w9873;
assign w9875 = w9859 & ~w9873;
assign w9876 = ~w9874 & ~w9875;
assign w9877 = ~w9845 & ~w9876;
assign w9878 = w9845 & w9876;
assign w9879 = ~w9877 & ~w9878;
assign w9880 = ~w9843 & w9879;
assign w9881 = w9843 & ~w9879;
assign w9882 = ~w9880 & ~w9881;
assign w9883 = ~w9807 & ~w9882;
assign w9884 = w9807 & w9882;
assign w9885 = ~w9883 & ~w9884;
assign w9886 = ~w9805 & w9885;
assign w9887 = w9805 & ~w9885;
assign w9888 = ~w9886 & ~w9887;
assign w9889 = ~w9725 & ~w9888;
assign w9890 = w9725 & w9888;
assign w9891 = ~w9889 & ~w9890;
assign w9892 = ~w1157 & ~w1546;
assign w9893 = ~w1547 & ~w9892;
assign w9894 = ~w1151 & ~w1154;
assign w9895 = ~w1155 & ~w9894;
assign w9896 = ~w1146 & ~w1148;
assign w9897 = ~w1149 & ~w9896;
assign w9898 = (w1130 & w1133) | (w1130 & w13574) | (w1133 & w13574);
assign w9899 = ~w1144 & ~w9898;
assign w9900 = ~w1047 & ~w1061;
assign w9901 = ~w1058 & ~w9900;
assign w9902 = ~w1080 & ~w1094;
assign w9903 = ~w1091 & ~w9902;
assign w9904 = ~w9901 & w9903;
assign w9905 = w9901 & ~w9903;
assign w9906 = ~w9904 & ~w9905;
assign w9907 = ~w9899 & ~w9906;
assign w9908 = ~w1144 & ~w9904;
assign w9909 = ~w9905 & w9908;
assign w9910 = ~w9898 & w9909;
assign w9911 = ~w9907 & ~w9910;
assign w9912 = (w1109 & w1112) | (w1109 & w13575) | (w1112 & w13575);
assign w9913 = ~w1119 & ~w9912;
assign w9914 = ~w978 & ~w992;
assign w9915 = ~w989 & ~w9914;
assign w9916 = ~w1011 & ~w1025;
assign w9917 = ~w1022 & ~w9916;
assign w9918 = ~w9915 & w9917;
assign w9919 = w9915 & ~w9917;
assign w9920 = ~w9918 & ~w9919;
assign w9921 = ~w9913 & ~w9920;
assign w9922 = ~w1119 & ~w9918;
assign w9923 = ~w9919 & w9922;
assign w9924 = ~w9912 & w9923;
assign w9925 = ~w9921 & ~w9924;
assign w9926 = ~w9911 & w9925;
assign w9927 = w9911 & ~w9925;
assign w9928 = ~w9926 & ~w9927;
assign w9929 = ~w9897 & ~w9928;
assign w9930 = w9897 & w9928;
assign w9931 = ~w9929 & ~w9930;
assign w9932 = ~w859 & ~w952;
assign w9933 = ~w953 & ~w9932;
assign w9934 = (w810 & w846) | (w810 & w13576) | (w846 & w13576);
assign w9935 = ~w857 & ~w9934;
assign w9936 = ~w839 & ~w843;
assign w9937 = ~w836 & ~w9936;
assign w9938 = ~w802 & ~w805;
assign w9939 = ~w808 & ~w9938;
assign w9940 = ~w9937 & w9939;
assign w9941 = w9937 & ~w9939;
assign w9942 = ~w9940 & ~w9941;
assign w9943 = ~w9935 & ~w9942;
assign w9944 = ~w857 & ~w9940;
assign w9945 = ~w9941 & w9944;
assign w9946 = ~w9934 & w9945;
assign w9947 = ~w9943 & ~w9946;
assign w9948 = (w892 & w928) | (w892 & w13577) | (w928 & w13577);
assign w9949 = ~w935 & ~w9948;
assign w9950 = ~w921 & ~w925;
assign w9951 = ~w918 & ~w9950;
assign w9952 = ~w884 & ~w887;
assign w9953 = ~w890 & ~w9952;
assign w9954 = ~w9951 & w9953;
assign w9955 = w9951 & ~w9953;
assign w9956 = ~w9954 & ~w9955;
assign w9957 = ~w9949 & ~w9956;
assign w9958 = ~w935 & ~w9954;
assign w9959 = ~w9955 & w9958;
assign w9960 = ~w9948 & w9959;
assign w9961 = ~w9957 & ~w9960;
assign w9962 = ~w9947 & w9961;
assign w9963 = w9947 & ~w9961;
assign w9964 = ~w9962 & ~w9963;
assign w9965 = ~w9933 & ~w9964;
assign w9966 = w9933 & w9964;
assign w9967 = ~w9965 & ~w9966;
assign w9968 = ~w9931 & w9967;
assign w9969 = w9931 & ~w9967;
assign w9970 = ~w9968 & ~w9969;
assign w9971 = ~w9895 & ~w9970;
assign w9972 = w9895 & w9970;
assign w9973 = ~w9971 & ~w9972;
assign w9974 = ~w1339 & ~w1529;
assign w9975 = ~w1531 & ~w9974;
assign w9976 = ~w1334 & ~w1336;
assign w9977 = ~w1337 & ~w9976;
assign w9978 = (w1318 & w1321) | (w1318 & w13578) | (w1321 & w13578);
assign w9979 = ~w1332 & ~w9978;
assign w9980 = ~w1260 & ~w1274;
assign w9981 = ~w1271 & ~w9980;
assign w9982 = ~w1293 & ~w1307;
assign w9983 = ~w1304 & ~w9982;
assign w9984 = ~w9981 & w9983;
assign w9985 = w9981 & ~w9983;
assign w9986 = ~w9984 & ~w9985;
assign w9987 = ~w9979 & ~w9986;
assign w9988 = ~w1332 & ~w9984;
assign w9989 = ~w9985 & w9988;
assign w9990 = ~w9978 & w9989;
assign w9991 = ~w9987 & ~w9990;
assign w9992 = (w1190 & w1226) | (w1190 & w13579) | (w1226 & w13579);
assign w9993 = ~w1233 & ~w9992;
assign w9994 = ~w1219 & ~w1223;
assign w9995 = ~w1216 & ~w9994;
assign w9996 = ~w1182 & ~w1185;
assign w9997 = ~w1188 & ~w9996;
assign w9998 = ~w9995 & w9997;
assign w9999 = w9995 & ~w9997;
assign w10000 = ~w9998 & ~w9999;
assign w10001 = ~w9993 & ~w10000;
assign w10002 = ~w1233 & ~w9998;
assign w10003 = ~w9999 & w10002;
assign w10004 = ~w9992 & w10003;
assign w10005 = ~w10001 & ~w10004;
assign w10006 = ~w9991 & w10005;
assign w10007 = w9991 & ~w10005;
assign w10008 = ~w10006 & ~w10007;
assign w10009 = ~w9977 & ~w10008;
assign w10010 = w9977 & w10008;
assign w10011 = ~w10009 & ~w10010;
assign w10012 = ~w1421 & ~w1514;
assign w10013 = ~w1515 & ~w10012;
assign w10014 = (w1372 & w1408) | (w1372 & w13580) | (w1408 & w13580);
assign w10015 = ~w1419 & ~w10014;
assign w10016 = ~w1401 & ~w1405;
assign w10017 = ~w1398 & ~w10016;
assign w10018 = ~w1364 & ~w1367;
assign w10019 = ~w1370 & ~w10018;
assign w10020 = ~w10017 & w10019;
assign w10021 = w10017 & ~w10019;
assign w10022 = ~w10020 & ~w10021;
assign w10023 = ~w10015 & ~w10022;
assign w10024 = ~w1419 & ~w10020;
assign w10025 = ~w10021 & w10024;
assign w10026 = ~w10014 & w10025;
assign w10027 = ~w10023 & ~w10026;
assign w10028 = (w1454 & w1490) | (w1454 & w13581) | (w1490 & w13581);
assign w10029 = ~w1497 & ~w10028;
assign w10030 = ~w1483 & ~w1487;
assign w10031 = ~w1480 & ~w10030;
assign w10032 = ~w1446 & ~w1449;
assign w10033 = ~w1452 & ~w10032;
assign w10034 = ~w10031 & w10033;
assign w10035 = w10031 & ~w10033;
assign w10036 = ~w10034 & ~w10035;
assign w10037 = ~w10029 & ~w10036;
assign w10038 = ~w1497 & ~w10034;
assign w10039 = ~w10035 & w10038;
assign w10040 = ~w10028 & w10039;
assign w10041 = ~w10037 & ~w10040;
assign w10042 = ~w10027 & w10041;
assign w10043 = w10027 & ~w10041;
assign w10044 = ~w10042 & ~w10043;
assign w10045 = ~w10013 & ~w10044;
assign w10046 = w10013 & w10044;
assign w10047 = ~w10045 & ~w10046;
assign w10048 = ~w10011 & w10047;
assign w10049 = w10011 & ~w10047;
assign w10050 = ~w10048 & ~w10049;
assign w10051 = ~w9975 & ~w10050;
assign w10052 = w9975 & w10050;
assign w10053 = ~w10051 & ~w10052;
assign w10054 = ~w9973 & w10053;
assign w10055 = w9973 & ~w10053;
assign w10056 = ~w10054 & ~w10055;
assign w10057 = ~w9893 & ~w10056;
assign w10058 = w9893 & w10056;
assign w10059 = ~w10057 & ~w10058;
assign w10060 = ~w9891 & w10059;
assign w10061 = w9891 & ~w10059;
assign w10062 = ~w10060 & ~w10061;
assign w10063 = ~w9723 & ~w10062;
assign w10064 = w9723 & w10062;
assign w10065 = ~w10063 & ~w10064;
assign w10066 = ~w9721 & w10065;
assign w10067 = w9721 & ~w10065;
assign w10068 = ~w10066 & ~w10067;
assign w10069 = ~w9377 & ~w10068;
assign w10070 = w9377 & w10068;
assign w10071 = ~w10069 & ~w10070;
assign w10072 = (~w8254 & w9375) | (~w8254 & w13888) | (w9375 & w13888);
assign w10073 = (w10071 & w9372) | (w10071 & w14065) | (w9372 & w14065);
assign w10074 = ~w9374 & w10073;
assign w10075 = ~w10072 & ~w10074;
assign w10076 = (~w8256 & w9369) | (~w8256 & w13889) | (w9369 & w13889);
assign w10077 = w8673 & w9369;
assign w10078 = ~w10076 & ~w10077;
assign w10079 = ~w9019 & ~w9363;
assign w10080 = ~w8675 & ~w10079;
assign w10081 = w9019 & w9363;
assign w10082 = ~w10080 & ~w10081;
assign w10083 = ~w9189 & ~w9357;
assign w10084 = ~w9021 & ~w10083;
assign w10085 = w9189 & w9357;
assign w10086 = ~w10084 & ~w10085;
assign w10087 = ~w9271 & ~w9351;
assign w10088 = ~w9191 & ~w10087;
assign w10089 = w9271 & w9351;
assign w10090 = ~w10088 & ~w10089;
assign w10091 = ~w9309 & ~w9345;
assign w10092 = ~w9273 & ~w10091;
assign w10093 = w9309 & w9345;
assign w10094 = ~w10092 & ~w10093;
assign w10095 = ~w9325 & ~w9339;
assign w10096 = ~w9311 & ~w10095;
assign w10097 = ~w9324 & ~w9338;
assign w10098 = w10097 & w12900;
assign w10099 = (~w10098 & w9311) | (~w10098 & w13049) | (w9311 & w13049);
assign w10100 = ~w8133 & ~w9329;
assign w10101 = ~w9326 & w10100;
assign w10102 = w9331 & ~w10101;
assign w10103 = (w9329 & w9326) | (w9329 & w13050) | (w9326 & w13050);
assign w10104 = ~w10102 & ~w10103;
assign w10105 = ~w8055 & ~w9315;
assign w10106 = ~w9312 & w10105;
assign w10107 = w9317 & ~w10106;
assign w10108 = (w9315 & w9312) | (w9315 & w13051) | (w9312 & w13051);
assign w10109 = ~w10107 & ~w10108;
assign w10110 = ~w10104 & w10109;
assign w10111 = w10104 & ~w10109;
assign w10112 = ~w10110 & ~w10111;
assign w10113 = ~w10099 & ~w10112;
assign w10114 = ~w10098 & ~w10110;
assign w10115 = ~w10111 & w10114;
assign w10116 = ~w10096 & w10115;
assign w10117 = ~w10113 & ~w10116;
assign w10118 = ~w9289 & ~w9303;
assign w10119 = (~w10118 & w9274) | (~w10118 & w12901) | (w9274 & w12901);
assign w10120 = ~w9288 & ~w9302;
assign w10121 = w10120 & w12902;
assign w10122 = (~w12901 & w13052) | (~w12901 & w13053) | (w13052 & w13053);
assign w10123 = ~w7869 & ~w9293;
assign w10124 = ~w9290 & w10123;
assign w10125 = w9295 & ~w10124;
assign w10126 = (w9293 & w9290) | (w9293 & w13054) | (w9290 & w13054);
assign w10127 = ~w10125 & ~w10126;
assign w10128 = ~w7968 & ~w9279;
assign w10129 = ~w9276 & w10128;
assign w10130 = w9281 & ~w10129;
assign w10131 = (w9279 & w9276) | (w9279 & w13055) | (w9276 & w13055);
assign w10132 = ~w10130 & ~w10131;
assign w10133 = ~w10127 & w10132;
assign w10134 = w10127 & ~w10132;
assign w10135 = ~w10133 & ~w10134;
assign w10136 = ~w10122 & ~w10135;
assign w10137 = ~w10121 & ~w10133;
assign w10138 = ~w10134 & w10137;
assign w10139 = ~w10119 & w10138;
assign w10140 = ~w10136 & ~w10139;
assign w10141 = ~w10117 & w10140;
assign w10142 = w10117 & ~w10140;
assign w10143 = ~w10141 & ~w10142;
assign w10144 = ~w10094 & ~w10143;
assign w10145 = w10094 & w10143;
assign w10146 = ~w10144 & ~w10145;
assign w10147 = ~w9229 & ~w9265;
assign w10148 = w9229 & w9265;
assign w10149 = (~w10148 & w9193) | (~w10148 & w12903) | (w9193 & w12903);
assign w10150 = ~w9245 & ~w9259;
assign w10151 = (~w10150 & w9230) | (~w10150 & w12904) | (w9230 & w12904);
assign w10152 = ~w9244 & ~w9258;
assign w10153 = w10152 & w12905;
assign w10154 = (~w12904 & w13056) | (~w12904 & w13057) | (w13056 & w13057);
assign w10155 = ~w7570 & ~w9249;
assign w10156 = ~w9246 & w10155;
assign w10157 = w9251 & ~w10156;
assign w10158 = (w9249 & w9246) | (w9249 & w13058) | (w9246 & w13058);
assign w10159 = ~w10157 & ~w10158;
assign w10160 = ~w7492 & ~w9235;
assign w10161 = ~w9232 & w10160;
assign w10162 = w9237 & ~w10161;
assign w10163 = (w9235 & w9232) | (w9235 & w13059) | (w9232 & w13059);
assign w10164 = ~w10162 & ~w10163;
assign w10165 = ~w10159 & w10164;
assign w10166 = w10159 & ~w10164;
assign w10167 = ~w10165 & ~w10166;
assign w10168 = ~w10154 & ~w10167;
assign w10169 = ~w10153 & ~w10165;
assign w10170 = ~w10166 & w10169;
assign w10171 = ~w10151 & w10170;
assign w10172 = ~w10168 & ~w10171;
assign w10173 = ~w9209 & ~w9223;
assign w10174 = (~w10173 & w9194) | (~w10173 & w12906) | (w9194 & w12906);
assign w10175 = ~w9208 & ~w9222;
assign w10176 = w10175 & w12907;
assign w10177 = (~w12906 & w13060) | (~w12906 & w13061) | (w13060 & w13061);
assign w10178 = ~w7754 & ~w9213;
assign w10179 = ~w9210 & w10178;
assign w10180 = w9215 & ~w10179;
assign w10181 = (w9213 & w9210) | (w9213 & w13062) | (w9210 & w13062);
assign w10182 = ~w10180 & ~w10181;
assign w10183 = ~w7779 & ~w9199;
assign w10184 = ~w9196 & w10183;
assign w10185 = w9201 & ~w10184;
assign w10186 = (w9199 & w9196) | (w9199 & w13063) | (w9196 & w13063);
assign w10187 = ~w10185 & ~w10186;
assign w10188 = ~w10182 & w10187;
assign w10189 = w10182 & ~w10187;
assign w10190 = ~w10188 & ~w10189;
assign w10191 = ~w10177 & ~w10190;
assign w10192 = ~w10176 & ~w10188;
assign w10193 = ~w10189 & w10192;
assign w10194 = ~w10174 & w10193;
assign w10195 = ~w10191 & ~w10194;
assign w10196 = ~w10172 & w10195;
assign w10197 = w10172 & ~w10195;
assign w10198 = ~w10196 & ~w10197;
assign w10199 = ~w10149 & ~w10198;
assign w10200 = w10149 & w10198;
assign w10201 = ~w10199 & ~w10200;
assign w10202 = ~w10146 & w10201;
assign w10203 = w10146 & ~w10201;
assign w10204 = ~w10202 & ~w10203;
assign w10205 = ~w10090 & ~w10204;
assign w10206 = w10090 & w10204;
assign w10207 = ~w10205 & ~w10206;
assign w10208 = ~w9103 & ~w9183;
assign w10209 = w9103 & w9183;
assign w10210 = (~w10209 & w9023) | (~w10209 & w12908) | (w9023 & w12908);
assign w10211 = ~w9141 & ~w9177;
assign w10212 = w9141 & w9177;
assign w10213 = (~w10212 & w9105) | (~w10212 & w12909) | (w9105 & w12909);
assign w10214 = ~w9157 & ~w9171;
assign w10215 = (~w10214 & w9142) | (~w10214 & w12910) | (w9142 & w12910);
assign w10216 = ~w9156 & ~w9170;
assign w10217 = w10216 & w12911;
assign w10218 = (~w12910 & w13064) | (~w12910 & w13065) | (w13064 & w13065);
assign w10219 = ~w6973 & ~w9161;
assign w10220 = ~w9158 & w10219;
assign w10221 = w9163 & ~w10220;
assign w10222 = (w9161 & w9158) | (w9161 & w13066) | (w9158 & w13066);
assign w10223 = ~w10221 & ~w10222;
assign w10224 = ~w6895 & ~w9147;
assign w10225 = ~w9144 & w10224;
assign w10226 = w9149 & ~w10225;
assign w10227 = (w9147 & w9144) | (w9147 & w13067) | (w9144 & w13067);
assign w10228 = ~w10226 & ~w10227;
assign w10229 = ~w10223 & w10228;
assign w10230 = w10223 & ~w10228;
assign w10231 = ~w10229 & ~w10230;
assign w10232 = ~w10218 & ~w10231;
assign w10233 = ~w10217 & ~w10229;
assign w10234 = ~w10230 & w10233;
assign w10235 = ~w10215 & w10234;
assign w10236 = ~w10232 & ~w10235;
assign w10237 = ~w9121 & ~w9135;
assign w10238 = (~w10237 & w9106) | (~w10237 & w12912) | (w9106 & w12912);
assign w10239 = ~w9120 & ~w9134;
assign w10240 = w10239 & w12913;
assign w10241 = (~w12912 & w13068) | (~w12912 & w13069) | (w13068 & w13069);
assign w10242 = ~w6708 & ~w9125;
assign w10243 = ~w9122 & w10242;
assign w10244 = w9127 & ~w10243;
assign w10245 = (w9125 & w9122) | (w9125 & w13070) | (w9122 & w13070);
assign w10246 = ~w10244 & ~w10245;
assign w10247 = ~w6807 & ~w9111;
assign w10248 = ~w9108 & w10247;
assign w10249 = w9113 & ~w10248;
assign w10250 = (w9111 & w9108) | (w9111 & w13071) | (w9108 & w13071);
assign w10251 = ~w10249 & ~w10250;
assign w10252 = ~w10246 & w10251;
assign w10253 = w10246 & ~w10251;
assign w10254 = ~w10252 & ~w10253;
assign w10255 = ~w10241 & ~w10254;
assign w10256 = ~w10240 & ~w10252;
assign w10257 = ~w10253 & w10256;
assign w10258 = ~w10238 & w10257;
assign w10259 = ~w10255 & ~w10258;
assign w10260 = ~w10236 & w10259;
assign w10261 = w10236 & ~w10259;
assign w10262 = ~w10260 & ~w10261;
assign w10263 = ~w10213 & ~w10262;
assign w10264 = w10213 & w10262;
assign w10265 = ~w10263 & ~w10264;
assign w10266 = ~w9061 & ~w9097;
assign w10267 = w9061 & w9097;
assign w10268 = (~w10267 & w9025) | (~w10267 & w12914) | (w9025 & w12914);
assign w10269 = ~w9077 & ~w9091;
assign w10270 = (~w10269 & w9062) | (~w10269 & w12915) | (w9062 & w12915);
assign w10271 = ~w9076 & ~w9090;
assign w10272 = w10271 & w12916;
assign w10273 = (~w12915 & w13072) | (~w12915 & w13073) | (w13072 & w13073);
assign w10274 = ~w7336 & ~w9081;
assign w10275 = ~w9078 & w10274;
assign w10276 = w9083 & ~w10275;
assign w10277 = (w9081 & w9078) | (w9081 & w13074) | (w9078 & w13074);
assign w10278 = ~w10276 & ~w10277;
assign w10279 = ~w7322 & ~w9067;
assign w10280 = ~w9064 & w10279;
assign w10281 = w9069 & ~w10280;
assign w10282 = (w9067 & w9064) | (w9067 & w13075) | (w9064 & w13075);
assign w10283 = ~w10281 & ~w10282;
assign w10284 = ~w10278 & w10283;
assign w10285 = w10278 & ~w10283;
assign w10286 = ~w10284 & ~w10285;
assign w10287 = ~w10273 & ~w10286;
assign w10288 = ~w10272 & ~w10284;
assign w10289 = ~w10285 & w10288;
assign w10290 = ~w10270 & w10289;
assign w10291 = ~w10287 & ~w10290;
assign w10292 = ~w9041 & ~w9055;
assign w10293 = (~w10292 & w9026) | (~w10292 & w12917) | (w9026 & w12917);
assign w10294 = ~w9040 & ~w9054;
assign w10295 = w10294 & w12918;
assign w10296 = (~w12917 & w13076) | (~w12917 & w13077) | (w13076 & w13077);
assign w10297 = ~w7366 & ~w9045;
assign w10298 = ~w9042 & w10297;
assign w10299 = w9047 & ~w10298;
assign w10300 = (w9045 & w9042) | (w9045 & w13078) | (w9042 & w13078);
assign w10301 = ~w10299 & ~w10300;
assign w10302 = ~w7391 & ~w9031;
assign w10303 = ~w9028 & w10302;
assign w10304 = w9033 & ~w10303;
assign w10305 = (w9031 & w9028) | (w9031 & w13079) | (w9028 & w13079);
assign w10306 = ~w10304 & ~w10305;
assign w10307 = ~w10301 & w10306;
assign w10308 = w10301 & ~w10306;
assign w10309 = ~w10307 & ~w10308;
assign w10310 = ~w10296 & ~w10309;
assign w10311 = ~w10295 & ~w10307;
assign w10312 = ~w10308 & w10311;
assign w10313 = ~w10293 & w10312;
assign w10314 = ~w10310 & ~w10313;
assign w10315 = ~w10291 & w10314;
assign w10316 = w10291 & ~w10314;
assign w10317 = ~w10315 & ~w10316;
assign w10318 = ~w10268 & ~w10317;
assign w10319 = w10268 & w10317;
assign w10320 = ~w10318 & ~w10319;
assign w10321 = ~w10265 & w10320;
assign w10322 = w10265 & ~w10320;
assign w10323 = ~w10321 & ~w10322;
assign w10324 = ~w10210 & ~w10323;
assign w10325 = w10210 & w10323;
assign w10326 = ~w10324 & ~w10325;
assign w10327 = ~w10207 & w10326;
assign w10328 = w10207 & ~w10326;
assign w10329 = ~w10327 & ~w10328;
assign w10330 = ~w10086 & ~w10329;
assign w10331 = w10086 & w10329;
assign w10332 = ~w10330 & ~w10331;
assign w10333 = ~w8845 & ~w9013;
assign w10334 = w8845 & w9013;
assign w10335 = (~w10334 & w8677) | (~w10334 & w12919) | (w8677 & w12919);
assign w10336 = ~w8927 & ~w9007;
assign w10337 = w8927 & w9007;
assign w10338 = (~w10337 & w8847) | (~w10337 & w12920) | (w8847 & w12920);
assign w10339 = ~w8965 & ~w9001;
assign w10340 = w8965 & w9001;
assign w10341 = (~w10340 & w8929) | (~w10340 & w12921) | (w8929 & w12921);
assign w10342 = ~w8981 & ~w8995;
assign w10343 = (~w10342 & w8966) | (~w10342 & w12922) | (w8966 & w12922);
assign w10344 = ~w8980 & ~w8994;
assign w10345 = w10344 & w12923;
assign w10346 = (~w12922 & w13080) | (~w12922 & w13081) | (w13080 & w13081);
assign w10347 = ~w5778 & ~w8985;
assign w10348 = ~w8982 & w10347;
assign w10349 = w8987 & ~w10348;
assign w10350 = (w8985 & w8982) | (w8985 & w13082) | (w8982 & w13082);
assign w10351 = ~w10349 & ~w10350;
assign w10352 = ~w5700 & ~w8971;
assign w10353 = ~w8968 & w10352;
assign w10354 = w8973 & ~w10353;
assign w10355 = (w8971 & w8968) | (w8971 & w13083) | (w8968 & w13083);
assign w10356 = ~w10354 & ~w10355;
assign w10357 = ~w10351 & w10356;
assign w10358 = w10351 & ~w10356;
assign w10359 = ~w10357 & ~w10358;
assign w10360 = ~w10346 & ~w10359;
assign w10361 = ~w10345 & ~w10357;
assign w10362 = ~w10358 & w10361;
assign w10363 = ~w10343 & w10362;
assign w10364 = ~w10360 & ~w10363;
assign w10365 = ~w8945 & ~w8959;
assign w10366 = (~w10365 & w8930) | (~w10365 & w12924) | (w8930 & w12924);
assign w10367 = ~w8944 & ~w8958;
assign w10368 = w10367 & w12925;
assign w10369 = (~w12924 & w13084) | (~w12924 & w13085) | (w13084 & w13085);
assign w10370 = ~w5513 & ~w8949;
assign w10371 = ~w8946 & w10370;
assign w10372 = w8951 & ~w10371;
assign w10373 = (w8949 & w8946) | (w8949 & w13086) | (w8946 & w13086);
assign w10374 = ~w10372 & ~w10373;
assign w10375 = ~w5612 & ~w8935;
assign w10376 = ~w8932 & w10375;
assign w10377 = w8937 & ~w10376;
assign w10378 = (w8935 & w8932) | (w8935 & w13087) | (w8932 & w13087);
assign w10379 = ~w10377 & ~w10378;
assign w10380 = ~w10374 & w10379;
assign w10381 = w10374 & ~w10379;
assign w10382 = ~w10380 & ~w10381;
assign w10383 = ~w10369 & ~w10382;
assign w10384 = ~w10368 & ~w10380;
assign w10385 = ~w10381 & w10384;
assign w10386 = ~w10366 & w10385;
assign w10387 = ~w10383 & ~w10386;
assign w10388 = ~w10364 & w10387;
assign w10389 = w10364 & ~w10387;
assign w10390 = ~w10388 & ~w10389;
assign w10391 = ~w10341 & ~w10390;
assign w10392 = w10341 & w10390;
assign w10393 = ~w10391 & ~w10392;
assign w10394 = ~w8885 & ~w8921;
assign w10395 = w8885 & w8921;
assign w10396 = (~w10395 & w8849) | (~w10395 & w12926) | (w8849 & w12926);
assign w10397 = ~w8901 & ~w8915;
assign w10398 = (~w10397 & w8886) | (~w10397 & w12927) | (w8886 & w12927);
assign w10399 = ~w8900 & ~w8914;
assign w10400 = w10399 & w12928;
assign w10401 = (~w12927 & w13088) | (~w12927 & w13089) | (w13088 & w13089);
assign w10402 = ~w5214 & ~w8905;
assign w10403 = ~w8902 & w10402;
assign w10404 = w8907 & ~w10403;
assign w10405 = (w8905 & w8902) | (w8905 & w13090) | (w8902 & w13090);
assign w10406 = ~w10404 & ~w10405;
assign w10407 = ~w5136 & ~w8891;
assign w10408 = ~w8888 & w10407;
assign w10409 = w8893 & ~w10408;
assign w10410 = (w8891 & w8888) | (w8891 & w13091) | (w8888 & w13091);
assign w10411 = ~w10409 & ~w10410;
assign w10412 = ~w10406 & w10411;
assign w10413 = w10406 & ~w10411;
assign w10414 = ~w10412 & ~w10413;
assign w10415 = ~w10401 & ~w10414;
assign w10416 = ~w10400 & ~w10412;
assign w10417 = ~w10413 & w10416;
assign w10418 = ~w10398 & w10417;
assign w10419 = ~w10415 & ~w10418;
assign w10420 = ~w8865 & ~w8879;
assign w10421 = (~w10420 & w8850) | (~w10420 & w12929) | (w8850 & w12929);
assign w10422 = ~w8864 & ~w8878;
assign w10423 = w10422 & w12930;
assign w10424 = (~w12929 & w13092) | (~w12929 & w13093) | (w13092 & w13093);
assign w10425 = ~w5398 & ~w8869;
assign w10426 = ~w8866 & w10425;
assign w10427 = w8871 & ~w10426;
assign w10428 = (w8869 & w8866) | (w8869 & w13094) | (w8866 & w13094);
assign w10429 = ~w10427 & ~w10428;
assign w10430 = ~w5423 & ~w8855;
assign w10431 = ~w8852 & w10430;
assign w10432 = w8857 & ~w10431;
assign w10433 = (w8855 & w8852) | (w8855 & w13095) | (w8852 & w13095);
assign w10434 = ~w10432 & ~w10433;
assign w10435 = ~w10429 & w10434;
assign w10436 = w10429 & ~w10434;
assign w10437 = ~w10435 & ~w10436;
assign w10438 = ~w10424 & ~w10437;
assign w10439 = ~w10423 & ~w10435;
assign w10440 = ~w10436 & w10439;
assign w10441 = ~w10421 & w10440;
assign w10442 = ~w10438 & ~w10441;
assign w10443 = ~w10419 & w10442;
assign w10444 = w10419 & ~w10442;
assign w10445 = ~w10443 & ~w10444;
assign w10446 = ~w10396 & ~w10445;
assign w10447 = w10396 & w10445;
assign w10448 = ~w10446 & ~w10447;
assign w10449 = ~w10393 & w10448;
assign w10450 = w10393 & ~w10448;
assign w10451 = ~w10449 & ~w10450;
assign w10452 = ~w10338 & ~w10451;
assign w10453 = w10338 & w10451;
assign w10454 = ~w10452 & ~w10453;
assign w10455 = ~w8759 & ~w8839;
assign w10456 = w8759 & w8839;
assign w10457 = (~w10456 & w8679) | (~w10456 & w12931) | (w8679 & w12931);
assign w10458 = ~w8797 & ~w8833;
assign w10459 = w8797 & w8833;
assign w10460 = (~w10459 & w8761) | (~w10459 & w12932) | (w8761 & w12932);
assign w10461 = ~w8813 & ~w8827;
assign w10462 = (~w10461 & w8798) | (~w10461 & w12933) | (w8798 & w12933);
assign w10463 = ~w8812 & ~w8826;
assign w10464 = w10463 & w12934;
assign w10465 = (~w12933 & w13096) | (~w12933 & w13097) | (w13096 & w13097);
assign w10466 = ~w6491 & ~w8817;
assign w10467 = ~w8814 & w10466;
assign w10468 = w8819 & ~w10467;
assign w10469 = (w8817 & w8814) | (w8817 & w13098) | (w8814 & w13098);
assign w10470 = ~w10468 & ~w10469;
assign w10471 = ~w6477 & ~w8803;
assign w10472 = ~w8800 & w10471;
assign w10473 = w8805 & ~w10472;
assign w10474 = (w8803 & w8800) | (w8803 & w13099) | (w8800 & w13099);
assign w10475 = ~w10473 & ~w10474;
assign w10476 = ~w10470 & w10475;
assign w10477 = w10470 & ~w10475;
assign w10478 = ~w10476 & ~w10477;
assign w10479 = ~w10465 & ~w10478;
assign w10480 = ~w10464 & ~w10476;
assign w10481 = ~w10477 & w10480;
assign w10482 = ~w10462 & w10481;
assign w10483 = ~w10479 & ~w10482;
assign w10484 = ~w8777 & ~w8791;
assign w10485 = (~w10484 & w8762) | (~w10484 & w12935) | (w8762 & w12935);
assign w10486 = ~w8776 & ~w8790;
assign w10487 = w10486 & w12936;
assign w10488 = (~w12935 & w13100) | (~w12935 & w13101) | (w13100 & w13101);
assign w10489 = ~w6428 & ~w8781;
assign w10490 = ~w8778 & w10489;
assign w10491 = w8783 & ~w10490;
assign w10492 = (w8781 & w8778) | (w8781 & w13102) | (w8778 & w13102);
assign w10493 = ~w10491 & ~w10492;
assign w10494 = ~w6453 & ~w8767;
assign w10495 = ~w8764 & w10494;
assign w10496 = w8769 & ~w10495;
assign w10497 = (w8767 & w8764) | (w8767 & w13103) | (w8764 & w13103);
assign w10498 = ~w10496 & ~w10497;
assign w10499 = ~w10493 & w10498;
assign w10500 = w10493 & ~w10498;
assign w10501 = ~w10499 & ~w10500;
assign w10502 = ~w10488 & ~w10501;
assign w10503 = ~w10487 & ~w10499;
assign w10504 = ~w10500 & w10503;
assign w10505 = ~w10485 & w10504;
assign w10506 = ~w10502 & ~w10505;
assign w10507 = ~w10483 & w10506;
assign w10508 = w10483 & ~w10506;
assign w10509 = ~w10507 & ~w10508;
assign w10510 = ~w10460 & ~w10509;
assign w10511 = w10460 & w10509;
assign w10512 = ~w10510 & ~w10511;
assign w10513 = ~w8717 & ~w8753;
assign w10514 = w8717 & w8753;
assign w10515 = (~w10514 & w8681) | (~w10514 & w12937) | (w8681 & w12937);
assign w10516 = ~w8733 & ~w8747;
assign w10517 = (~w10516 & w8718) | (~w10516 & w12938) | (w8718 & w12938);
assign w10518 = ~w8732 & ~w8746;
assign w10519 = w10518 & w12939;
assign w10520 = (~w12938 & w13104) | (~w12938 & w13105) | (w13104 & w13105);
assign w10521 = ~w6550 & ~w8737;
assign w10522 = ~w8734 & w10521;
assign w10523 = w8739 & ~w10522;
assign w10524 = (w8737 & w8734) | (w8737 & w13106) | (w8734 & w13106);
assign w10525 = ~w10523 & ~w10524;
assign w10526 = ~w6536 & ~w8723;
assign w10527 = ~w8720 & w10526;
assign w10528 = w8725 & ~w10527;
assign w10529 = (w8723 & w8720) | (w8723 & w13107) | (w8720 & w13107);
assign w10530 = ~w10528 & ~w10529;
assign w10531 = ~w10525 & w10530;
assign w10532 = w10525 & ~w10530;
assign w10533 = ~w10531 & ~w10532;
assign w10534 = ~w10520 & ~w10533;
assign w10535 = ~w10519 & ~w10531;
assign w10536 = ~w10532 & w10535;
assign w10537 = ~w10517 & w10536;
assign w10538 = ~w10534 & ~w10537;
assign w10539 = ~w8697 & ~w8711;
assign w10540 = (~w10539 & w8682) | (~w10539 & w12940) | (w8682 & w12940);
assign w10541 = ~w8696 & ~w8710;
assign w10542 = w10541 & w12941;
assign w10543 = (~w12940 & w13108) | (~w12940 & w13109) | (w13108 & w13109);
assign w10544 = ~w6580 & ~w8701;
assign w10545 = ~w8698 & w10544;
assign w10546 = w8703 & ~w10545;
assign w10547 = (w8701 & w8698) | (w8701 & w13110) | (w8698 & w13110);
assign w10548 = ~w10546 & ~w10547;
assign w10549 = ~w6605 & ~w8687;
assign w10550 = ~w8684 & w10549;
assign w10551 = w8689 & ~w10550;
assign w10552 = (w8687 & w8684) | (w8687 & w13111) | (w8684 & w13111);
assign w10553 = ~w10551 & ~w10552;
assign w10554 = ~w10548 & w10553;
assign w10555 = w10548 & ~w10553;
assign w10556 = ~w10554 & ~w10555;
assign w10557 = ~w10543 & ~w10556;
assign w10558 = ~w10542 & ~w10554;
assign w10559 = ~w10555 & w10558;
assign w10560 = ~w10540 & w10559;
assign w10561 = ~w10557 & ~w10560;
assign w10562 = ~w10538 & w10561;
assign w10563 = w10538 & ~w10561;
assign w10564 = ~w10562 & ~w10563;
assign w10565 = ~w10515 & ~w10564;
assign w10566 = w10515 & w10564;
assign w10567 = ~w10565 & ~w10566;
assign w10568 = ~w10512 & w10567;
assign w10569 = w10512 & ~w10567;
assign w10570 = ~w10568 & ~w10569;
assign w10571 = ~w10457 & ~w10570;
assign w10572 = w10457 & w10570;
assign w10573 = ~w10571 & ~w10572;
assign w10574 = ~w10454 & w10573;
assign w10575 = w10454 & ~w10573;
assign w10576 = ~w10574 & ~w10575;
assign w10577 = ~w10335 & ~w10576;
assign w10578 = w10335 & w10576;
assign w10579 = ~w10577 & ~w10578;
assign w10580 = ~w10332 & w10579;
assign w10581 = w10332 & ~w10579;
assign w10582 = ~w10580 & ~w10581;
assign w10583 = ~w10082 & ~w10582;
assign w10584 = w10082 & w10582;
assign w10585 = ~w10583 & ~w10584;
assign w10586 = ~w8666 & ~w8669;
assign w10587 = ~w8258 & ~w10586;
assign w10588 = ~w8498 & w8666;
assign w10589 = ~w8497 & w10588;
assign w10590 = ~w10587 & ~w10589;
assign w10591 = ~w8491 & ~w8494;
assign w10592 = (w8491 & w8409) | (w8491 & w13890) | (w8409 & w13890);
assign w10593 = ~w8410 & w10592;
assign w10594 = (~w10593 & w10591) | (~w10593 & w13891) | (w10591 & w13891);
assign w10595 = ~w8326 & ~w8406;
assign w10596 = w8326 & w8406;
assign w10597 = (~w10596 & w8262) | (~w10596 & w12942) | (w8262 & w12942);
assign w10598 = ~w8364 & ~w8400;
assign w10599 = w8364 & w8400;
assign w10600 = (~w10599 & w8328) | (~w10599 & w12943) | (w8328 & w12943);
assign w10601 = ~w8380 & ~w8394;
assign w10602 = (~w10601 & w8365) | (~w10601 & w12944) | (w8365 & w12944);
assign w10603 = ~w8379 & ~w8393;
assign w10604 = w10603 & w12945;
assign w10605 = (~w12944 & w13112) | (~w12944 & w13113) | (w13112 & w13113);
assign w10606 = ~w4183 & ~w8384;
assign w10607 = ~w8381 & w10606;
assign w10608 = w8386 & ~w10607;
assign w10609 = (w8384 & w8381) | (w8384 & w13114) | (w8381 & w13114);
assign w10610 = ~w10608 & ~w10609;
assign w10611 = ~w4105 & ~w8370;
assign w10612 = ~w8367 & w10611;
assign w10613 = w8372 & ~w10612;
assign w10614 = (w8370 & w8367) | (w8370 & w13115) | (w8367 & w13115);
assign w10615 = ~w10613 & ~w10614;
assign w10616 = ~w10610 & w10615;
assign w10617 = w10610 & ~w10615;
assign w10618 = ~w10616 & ~w10617;
assign w10619 = ~w10605 & ~w10618;
assign w10620 = ~w10604 & ~w10616;
assign w10621 = ~w10617 & w10620;
assign w10622 = ~w10602 & w10621;
assign w10623 = ~w10619 & ~w10622;
assign w10624 = ~w8344 & ~w8358;
assign w10625 = (~w10624 & w8329) | (~w10624 & w12946) | (w8329 & w12946);
assign w10626 = ~w8343 & ~w8357;
assign w10627 = w10626 & w12947;
assign w10628 = (~w12946 & w13116) | (~w12946 & w13117) | (w13116 & w13117);
assign w10629 = ~w3918 & ~w8348;
assign w10630 = ~w8345 & w10629;
assign w10631 = w8350 & ~w10630;
assign w10632 = (w8348 & w8345) | (w8348 & w13118) | (w8345 & w13118);
assign w10633 = ~w10631 & ~w10632;
assign w10634 = ~w4017 & ~w8334;
assign w10635 = ~w8331 & w10634;
assign w10636 = w8336 & ~w10635;
assign w10637 = (w8334 & w8331) | (w8334 & w13119) | (w8331 & w13119);
assign w10638 = ~w10636 & ~w10637;
assign w10639 = ~w10633 & w10638;
assign w10640 = w10633 & ~w10638;
assign w10641 = ~w10639 & ~w10640;
assign w10642 = ~w10628 & ~w10641;
assign w10643 = ~w10627 & ~w10639;
assign w10644 = ~w10640 & w10643;
assign w10645 = ~w10625 & w10644;
assign w10646 = ~w10642 & ~w10645;
assign w10647 = ~w10623 & w10646;
assign w10648 = w10623 & ~w10646;
assign w10649 = ~w10647 & ~w10648;
assign w10650 = ~w10600 & ~w10649;
assign w10651 = w10600 & w10649;
assign w10652 = ~w10650 & ~w10651;
assign w10653 = ~w8284 & ~w8320;
assign w10654 = w8284 & ~w8318;
assign w10655 = ~w8319 & w10654;
assign w10656 = (~w10655 & w8264) | (~w10655 & w12948) | (w8264 & w12948);
assign w10657 = ~w3833 & w8278;
assign w10658 = (w8275 & ~w10657) | (w8275 & w12949) | (~w10657 & w12949);
assign w10659 = ~w8266 & ~w8278;
assign w10660 = ~w10658 & ~w10659;
assign w10661 = ~w8268 & ~w8270;
assign w10662 = ~w10660 & w10661;
assign w10663 = (w10657 & w13892) | (w10657 & w13893) | (w13892 & w13893);
assign w10664 = ~w10659 & w10663;
assign w10665 = ~w10662 & ~w10664;
assign w10666 = ~w8300 & ~w8314;
assign w10667 = ~w8286 & ~w10666;
assign w10668 = ~w8299 & ~w8313;
assign w10669 = w10668 & w12950;
assign w10670 = ~w3700 & ~w8304;
assign w10671 = ~w8301 & w10670;
assign w10672 = w8306 & ~w10671;
assign w10673 = (w8304 & w8301) | (w8304 & w13430) | (w8301 & w13430);
assign w10674 = ~w10672 & ~w10673;
assign w10675 = ~w3622 & ~w8290;
assign w10676 = ~w8287 & w10675;
assign w10677 = w8292 & ~w10676;
assign w10678 = (w8290 & w8287) | (w8290 & w13431) | (w8287 & w13431);
assign w10679 = ~w10677 & ~w10678;
assign w10680 = ~w10674 & w10679;
assign w10681 = w10674 & ~w10679;
assign w10682 = ~w10680 & ~w10681;
assign w10683 = (~w10682 & w10667) | (~w10682 & w12951) | (w10667 & w12951);
assign w10684 = ~w10669 & ~w10680;
assign w10685 = ~w10681 & w10684;
assign w10686 = ~w10667 & w10685;
assign w10687 = ~w10683 & ~w10686;
assign w10688 = ~w10665 & ~w10687;
assign w10689 = w10665 & w10687;
assign w10690 = ~w10688 & ~w10689;
assign w10691 = ~w10656 & w10690;
assign w10692 = w10656 & ~w10690;
assign w10693 = ~w10691 & ~w10692;
assign w10694 = ~w10652 & w10693;
assign w10695 = w10652 & ~w10693;
assign w10696 = ~w10694 & ~w10695;
assign w10697 = ~w10597 & ~w10696;
assign w10698 = w10597 & w10696;
assign w10699 = ~w10697 & ~w10698;
assign w10700 = ~w8449 & ~w8485;
assign w10701 = ~w8413 & ~w10700;
assign w10702 = w8449 & w8485;
assign w10703 = ~w10701 & ~w10702;
assign w10704 = ~w8465 & ~w8479;
assign w10705 = ~w8451 & ~w10704;
assign w10706 = ~w8464 & ~w8478;
assign w10707 = w10706 & w13894;
assign w10708 = ~w3320 & ~w8469;
assign w10709 = ~w8466 & w10708;
assign w10710 = w8471 & ~w10709;
assign w10711 = (w8469 & w8466) | (w8469 & w13895) | (w8466 & w13895);
assign w10712 = ~w10710 & ~w10711;
assign w10713 = ~w3242 & ~w8455;
assign w10714 = ~w8452 & w10713;
assign w10715 = w8457 & ~w10714;
assign w10716 = (w8455 & w8452) | (w8455 & w13896) | (w8452 & w13896);
assign w10717 = ~w10715 & ~w10716;
assign w10718 = ~w10712 & w10717;
assign w10719 = w10712 & ~w10717;
assign w10720 = ~w10718 & ~w10719;
assign w10721 = (~w10720 & w10705) | (~w10720 & w13897) | (w10705 & w13897);
assign w10722 = ~w10707 & ~w10718;
assign w10723 = ~w10719 & w10722;
assign w10724 = ~w10705 & w10723;
assign w10725 = ~w10721 & ~w10724;
assign w10726 = ~w8429 & ~w8443;
assign w10727 = ~w8415 & ~w10726;
assign w10728 = ~w8428 & ~w8442;
assign w10729 = w10728 & w13898;
assign w10730 = ~w3504 & ~w8433;
assign w10731 = ~w8430 & w10730;
assign w10732 = w8435 & ~w10731;
assign w10733 = (w8433 & w8430) | (w8433 & w13899) | (w8430 & w13899);
assign w10734 = ~w10732 & ~w10733;
assign w10735 = ~w3529 & ~w8419;
assign w10736 = ~w8416 & w10735;
assign w10737 = w8421 & ~w10736;
assign w10738 = (w8419 & w8416) | (w8419 & w13900) | (w8416 & w13900);
assign w10739 = ~w10737 & ~w10738;
assign w10740 = ~w10734 & w10739;
assign w10741 = w10734 & ~w10739;
assign w10742 = ~w10740 & ~w10741;
assign w10743 = (~w10742 & w10727) | (~w10742 & w13901) | (w10727 & w13901);
assign w10744 = ~w10729 & ~w10740;
assign w10745 = ~w10741 & w10744;
assign w10746 = ~w10727 & w10745;
assign w10747 = ~w10743 & ~w10746;
assign w10748 = ~w10725 & w10747;
assign w10749 = w10725 & ~w10747;
assign w10750 = ~w10748 & ~w10749;
assign w10751 = ~w10703 & ~w10750;
assign w10752 = w10703 & w10750;
assign w10753 = ~w10751 & ~w10752;
assign w10754 = ~w10699 & w10753;
assign w10755 = ~w10697 & ~w10753;
assign w10756 = ~w10698 & w10755;
assign w10757 = ~w10754 & ~w10756;
assign w10758 = ~w10594 & ~w10757;
assign w10759 = w10594 & w10757;
assign w10760 = ~w10758 & ~w10759;
assign w10761 = ~w8580 & ~w8660;
assign w10762 = ~w8500 & ~w10761;
assign w10763 = w8580 & w8660;
assign w10764 = ~w10762 & ~w10763;
assign w10765 = ~w8618 & ~w8654;
assign w10766 = ~w8582 & ~w10765;
assign w10767 = w8618 & w8654;
assign w10768 = ~w10766 & ~w10767;
assign w10769 = ~w8634 & ~w8648;
assign w10770 = ~w8620 & ~w10769;
assign w10771 = ~w8633 & ~w8647;
assign w10772 = w10771 & w13582;
assign w10773 = (~w10772 & w8620) | (~w10772 & w13902) | (w8620 & w13902);
assign w10774 = ~w4915 & ~w8638;
assign w10775 = ~w8635 & w10774;
assign w10776 = w8640 & ~w10775;
assign w10777 = (w8638 & w8635) | (w8638 & w13903) | (w8635 & w13903);
assign w10778 = ~w10776 & ~w10777;
assign w10779 = ~w4901 & ~w8624;
assign w10780 = ~w8621 & w10779;
assign w10781 = w8626 & ~w10780;
assign w10782 = (w8624 & w8621) | (w8624 & w13904) | (w8621 & w13904);
assign w10783 = ~w10781 & ~w10782;
assign w10784 = ~w10778 & w10783;
assign w10785 = w10778 & ~w10783;
assign w10786 = ~w10784 & ~w10785;
assign w10787 = ~w10773 & ~w10786;
assign w10788 = ~w10772 & ~w10784;
assign w10789 = ~w10785 & w10788;
assign w10790 = ~w10770 & w10789;
assign w10791 = ~w10787 & ~w10790;
assign w10792 = ~w8598 & ~w8612;
assign w10793 = (~w10792 & w8583) | (~w10792 & w13583) | (w8583 & w13583);
assign w10794 = ~w8597 & ~w8611;
assign w10795 = w10794 & w13584;
assign w10796 = ~w10795 & ~w10793;
assign w10797 = ~w4853 & ~w8602;
assign w10798 = ~w8599 & w10797;
assign w10799 = w8604 & ~w10798;
assign w10800 = (w8602 & w8599) | (w8602 & w13905) | (w8599 & w13905);
assign w10801 = ~w10799 & ~w10800;
assign w10802 = ~w4878 & ~w8588;
assign w10803 = ~w8585 & w10802;
assign w10804 = w8590 & ~w10803;
assign w10805 = (w8588 & w8585) | (w8588 & w13906) | (w8585 & w13906);
assign w10806 = ~w10804 & ~w10805;
assign w10807 = ~w10801 & w10806;
assign w10808 = w10801 & ~w10806;
assign w10809 = ~w10807 & ~w10808;
assign w10810 = ~w10796 & ~w10809;
assign w10811 = ~w10795 & ~w10807;
assign w10812 = ~w10808 & w10811;
assign w10813 = ~w10793 & w10812;
assign w10814 = ~w10810 & ~w10813;
assign w10815 = ~w10791 & w10814;
assign w10816 = w10791 & ~w10814;
assign w10817 = ~w10815 & ~w10816;
assign w10818 = ~w10768 & ~w10817;
assign w10819 = w10768 & w10817;
assign w10820 = ~w10818 & ~w10819;
assign w10821 = ~w8538 & ~w8574;
assign w10822 = w8538 & w8574;
assign w10823 = (~w10822 & w8502) | (~w10822 & w13907) | (w8502 & w13907);
assign w10824 = ~w8554 & ~w8568;
assign w10825 = ~w8540 & ~w10824;
assign w10826 = ~w8553 & ~w8567;
assign w10827 = w10826 & w13585;
assign w10828 = (~w10827 & w8540) | (~w10827 & w13908) | (w8540 & w13908);
assign w10829 = ~w4974 & ~w8558;
assign w10830 = ~w8555 & w10829;
assign w10831 = w8560 & ~w10830;
assign w10832 = (w8558 & w8555) | (w8558 & w13909) | (w8555 & w13909);
assign w10833 = ~w10831 & ~w10832;
assign w10834 = ~w4960 & ~w8544;
assign w10835 = ~w8541 & w10834;
assign w10836 = w8546 & ~w10835;
assign w10837 = (w8544 & w8541) | (w8544 & w13910) | (w8541 & w13910);
assign w10838 = ~w10836 & ~w10837;
assign w10839 = ~w10833 & w10838;
assign w10840 = w10833 & ~w10838;
assign w10841 = ~w10839 & ~w10840;
assign w10842 = ~w10828 & ~w10841;
assign w10843 = ~w10827 & ~w10839;
assign w10844 = ~w10840 & w10843;
assign w10845 = ~w10825 & w10844;
assign w10846 = ~w10842 & ~w10845;
assign w10847 = ~w8518 & ~w8532;
assign w10848 = (~w10847 & w8503) | (~w10847 & w13586) | (w8503 & w13586);
assign w10849 = ~w8517 & ~w8531;
assign w10850 = w10849 & w13587;
assign w10851 = ~w10850 & ~w10848;
assign w10852 = ~w5004 & ~w8522;
assign w10853 = ~w8519 & w10852;
assign w10854 = w8524 & ~w10853;
assign w10855 = (w8522 & w8519) | (w8522 & w13911) | (w8519 & w13911);
assign w10856 = ~w10854 & ~w10855;
assign w10857 = ~w5029 & ~w8508;
assign w10858 = ~w8505 & w10857;
assign w10859 = w8510 & ~w10858;
assign w10860 = (w8508 & w8505) | (w8508 & w13912) | (w8505 & w13912);
assign w10861 = ~w10859 & ~w10860;
assign w10862 = ~w10856 & w10861;
assign w10863 = w10856 & ~w10861;
assign w10864 = ~w10862 & ~w10863;
assign w10865 = ~w10851 & ~w10864;
assign w10866 = ~w10850 & ~w10862;
assign w10867 = ~w10863 & w10866;
assign w10868 = ~w10848 & w10867;
assign w10869 = ~w10865 & ~w10868;
assign w10870 = ~w10846 & w10869;
assign w10871 = w10846 & ~w10869;
assign w10872 = ~w10870 & ~w10871;
assign w10873 = ~w10823 & ~w10872;
assign w10874 = w10823 & w10872;
assign w10875 = ~w10873 & ~w10874;
assign w10876 = ~w10820 & w10875;
assign w10877 = w10820 & ~w10875;
assign w10878 = ~w10876 & ~w10877;
assign w10879 = ~w10764 & ~w10878;
assign w10880 = w10764 & w10878;
assign w10881 = ~w10879 & ~w10880;
assign w10882 = ~w10760 & w10881;
assign w10883 = (~w10881 & w10757) | (~w10881 & w13913) | (w10757 & w13913);
assign w10884 = ~w10759 & w10883;
assign w10885 = ~w10882 & ~w10884;
assign w10886 = ~w10590 & ~w10885;
assign w10887 = w10590 & w10885;
assign w10888 = ~w10886 & ~w10887;
assign w10889 = ~w10585 & w10888;
assign w10890 = w10585 & ~w10888;
assign w10891 = ~w10889 & ~w10890;
assign w10892 = ~w10078 & ~w10891;
assign w10893 = w10078 & w10891;
assign w10894 = ~w10892 & ~w10893;
assign w10895 = ~w9721 & ~w10065;
assign w10896 = ~w9377 & ~w10895;
assign w10897 = w9721 & w10065;
assign w10898 = ~w10896 & ~w10897;
assign w10899 = ~w9891 & ~w10059;
assign w10900 = ~w9723 & ~w10899;
assign w10901 = w9891 & w10059;
assign w10902 = ~w10900 & ~w10901;
assign w10903 = ~w9973 & ~w10053;
assign w10904 = ~w9893 & ~w10903;
assign w10905 = w9973 & w10053;
assign w10906 = ~w10904 & ~w10905;
assign w10907 = ~w10011 & ~w10047;
assign w10908 = ~w9975 & ~w10907;
assign w10909 = w10011 & w10047;
assign w10910 = ~w10908 & ~w10909;
assign w10911 = ~w10027 & ~w10041;
assign w10912 = ~w10013 & ~w10911;
assign w10913 = ~w10026 & ~w10040;
assign w10914 = w10913 & w13588;
assign w10915 = (~w10914 & w10013) | (~w10914 & w13737) | (w10013 & w13737);
assign w10916 = ~w1497 & ~w10031;
assign w10917 = ~w10028 & w10916;
assign w10918 = w10033 & ~w10917;
assign w10919 = (w10031 & w10028) | (w10031 & w13738) | (w10028 & w13738);
assign w10920 = ~w10918 & ~w10919;
assign w10921 = ~w1419 & ~w10017;
assign w10922 = ~w10014 & w10921;
assign w10923 = w10019 & ~w10922;
assign w10924 = (w10017 & w10014) | (w10017 & w13739) | (w10014 & w13739);
assign w10925 = ~w10923 & ~w10924;
assign w10926 = ~w10920 & w10925;
assign w10927 = w10920 & ~w10925;
assign w10928 = ~w10926 & ~w10927;
assign w10929 = ~w10915 & ~w10928;
assign w10930 = ~w10914 & ~w10926;
assign w10931 = ~w10927 & w10930;
assign w10932 = ~w10912 & w10931;
assign w10933 = ~w10929 & ~w10932;
assign w10934 = ~w9991 & ~w10005;
assign w10935 = (~w10934 & w9976) | (~w10934 & w13589) | (w9976 & w13589);
assign w10936 = ~w9990 & ~w10004;
assign w10937 = w10936 & w13590;
assign w10938 = ~w10937 & ~w10935;
assign w10939 = ~w1233 & ~w9995;
assign w10940 = ~w9992 & w10939;
assign w10941 = w9997 & ~w10940;
assign w10942 = (w9995 & w9992) | (w9995 & w13740) | (w9992 & w13740);
assign w10943 = ~w10941 & ~w10942;
assign w10944 = ~w1332 & ~w9981;
assign w10945 = ~w9978 & w10944;
assign w10946 = w9983 & ~w10945;
assign w10947 = (w9981 & w9978) | (w9981 & w13741) | (w9978 & w13741);
assign w10948 = ~w10946 & ~w10947;
assign w10949 = ~w10943 & w10948;
assign w10950 = w10943 & ~w10948;
assign w10951 = ~w10949 & ~w10950;
assign w10952 = ~w10938 & ~w10951;
assign w10953 = ~w10937 & ~w10949;
assign w10954 = ~w10950 & w10953;
assign w10955 = ~w10935 & w10954;
assign w10956 = ~w10952 & ~w10955;
assign w10957 = ~w10933 & w10956;
assign w10958 = w10933 & ~w10956;
assign w10959 = ~w10957 & ~w10958;
assign w10960 = ~w10910 & ~w10959;
assign w10961 = w10910 & w10959;
assign w10962 = ~w10960 & ~w10961;
assign w10963 = ~w9931 & ~w9967;
assign w10964 = ~w9895 & ~w10963;
assign w10965 = w9931 & w9967;
assign w10966 = ~w10964 & ~w10965;
assign w10967 = ~w9947 & ~w9961;
assign w10968 = ~w9933 & ~w10967;
assign w10969 = ~w9946 & ~w9960;
assign w10970 = w10969 & w13591;
assign w10971 = (~w10970 & w9933) | (~w10970 & w13742) | (w9933 & w13742);
assign w10972 = ~w935 & ~w9951;
assign w10973 = ~w9948 & w10972;
assign w10974 = w9953 & ~w10973;
assign w10975 = (w9951 & w9948) | (w9951 & w13743) | (w9948 & w13743);
assign w10976 = ~w10974 & ~w10975;
assign w10977 = ~w857 & ~w9937;
assign w10978 = ~w9934 & w10977;
assign w10979 = w9939 & ~w10978;
assign w10980 = (w9937 & w9934) | (w9937 & w13744) | (w9934 & w13744);
assign w10981 = ~w10979 & ~w10980;
assign w10982 = ~w10976 & w10981;
assign w10983 = w10976 & ~w10981;
assign w10984 = ~w10982 & ~w10983;
assign w10985 = ~w10971 & ~w10984;
assign w10986 = ~w10970 & ~w10982;
assign w10987 = ~w10983 & w10986;
assign w10988 = ~w10968 & w10987;
assign w10989 = ~w10985 & ~w10988;
assign w10990 = ~w9911 & ~w9925;
assign w10991 = (~w10990 & w9896) | (~w10990 & w13592) | (w9896 & w13592);
assign w10992 = ~w9910 & ~w9924;
assign w10993 = w10992 & w13593;
assign w10994 = ~w10993 & ~w10991;
assign w10995 = ~w1119 & ~w9915;
assign w10996 = ~w9912 & w10995;
assign w10997 = w9917 & ~w10996;
assign w10998 = (w9915 & w9912) | (w9915 & w13745) | (w9912 & w13745);
assign w10999 = ~w10997 & ~w10998;
assign w11000 = ~w1144 & ~w9901;
assign w11001 = ~w9898 & w11000;
assign w11002 = w9903 & ~w11001;
assign w11003 = (w9901 & w9898) | (w9901 & w13746) | (w9898 & w13746);
assign w11004 = ~w11002 & ~w11003;
assign w11005 = ~w10999 & w11004;
assign w11006 = w10999 & ~w11004;
assign w11007 = ~w11005 & ~w11006;
assign w11008 = ~w10994 & ~w11007;
assign w11009 = ~w10993 & ~w11005;
assign w11010 = ~w11006 & w11009;
assign w11011 = ~w10991 & w11010;
assign w11012 = ~w11008 & ~w11011;
assign w11013 = ~w10989 & w11012;
assign w11014 = w10989 & ~w11012;
assign w11015 = ~w11013 & ~w11014;
assign w11016 = ~w10966 & ~w11015;
assign w11017 = w10966 & w11015;
assign w11018 = ~w11016 & ~w11017;
assign w11019 = ~w10962 & w11018;
assign w11020 = w10962 & ~w11018;
assign w11021 = ~w11019 & ~w11020;
assign w11022 = ~w10906 & ~w11021;
assign w11023 = w10906 & w11021;
assign w11024 = ~w11022 & ~w11023;
assign w11025 = ~w9805 & ~w9885;
assign w11026 = ~w9725 & ~w11025;
assign w11027 = w9805 & w9885;
assign w11028 = ~w11026 & ~w11027;
assign w11029 = ~w9843 & ~w9879;
assign w11030 = ~w9807 & ~w11029;
assign w11031 = w9843 & w9879;
assign w11032 = ~w11030 & ~w11031;
assign w11033 = ~w9859 & ~w9873;
assign w11034 = ~w9845 & ~w11033;
assign w11035 = ~w9858 & ~w9872;
assign w11036 = w11035 & w13594;
assign w11037 = (~w11036 & w9845) | (~w11036 & w13747) | (w9845 & w13747);
assign w11038 = ~w339 & ~w9863;
assign w11039 = ~w9860 & w11038;
assign w11040 = w9865 & ~w11039;
assign w11041 = (w9863 & w9860) | (w9863 & w13748) | (w9860 & w13748);
assign w11042 = ~w11040 & ~w11041;
assign w11043 = ~w261 & ~w9849;
assign w11044 = ~w9846 & w11043;
assign w11045 = w9851 & ~w11044;
assign w11046 = (w9849 & w9846) | (w9849 & w13749) | (w9846 & w13749);
assign w11047 = ~w11045 & ~w11046;
assign w11048 = ~w11042 & w11047;
assign w11049 = w11042 & ~w11047;
assign w11050 = ~w11048 & ~w11049;
assign w11051 = ~w11037 & ~w11050;
assign w11052 = ~w11036 & ~w11048;
assign w11053 = ~w11049 & w11052;
assign w11054 = ~w11034 & w11053;
assign w11055 = ~w11051 & ~w11054;
assign w11056 = ~w9823 & ~w9837;
assign w11057 = (~w11056 & w9808) | (~w11056 & w13595) | (w9808 & w13595);
assign w11058 = ~w9822 & ~w9836;
assign w11059 = w11058 & w13596;
assign w11060 = ~w11059 & ~w11057;
assign w11061 = ~w75 & ~w9827;
assign w11062 = ~w9824 & w11061;
assign w11063 = w9829 & ~w11062;
assign w11064 = (w9827 & w9824) | (w9827 & w13750) | (w9824 & w13750);
assign w11065 = ~w11063 & ~w11064;
assign w11066 = ~w174 & ~w9813;
assign w11067 = ~w9810 & w11066;
assign w11068 = w9815 & ~w11067;
assign w11069 = (w9813 & w9810) | (w9813 & w13751) | (w9810 & w13751);
assign w11070 = ~w11068 & ~w11069;
assign w11071 = ~w11065 & w11070;
assign w11072 = w11065 & ~w11070;
assign w11073 = ~w11071 & ~w11072;
assign w11074 = ~w11060 & ~w11073;
assign w11075 = ~w11059 & ~w11071;
assign w11076 = ~w11072 & w11075;
assign w11077 = ~w11057 & w11076;
assign w11078 = ~w11074 & ~w11077;
assign w11079 = ~w11055 & w11078;
assign w11080 = w11055 & ~w11078;
assign w11081 = ~w11079 & ~w11080;
assign w11082 = ~w11032 & ~w11081;
assign w11083 = w11032 & w11081;
assign w11084 = ~w11082 & ~w11083;
assign w11085 = ~w9763 & ~w9799;
assign w11086 = ~w9727 & ~w11085;
assign w11087 = w9763 & w9799;
assign w11088 = ~w11086 & ~w11087;
assign w11089 = ~w9779 & ~w9793;
assign w11090 = ~w9765 & ~w11089;
assign w11091 = ~w9778 & ~w9792;
assign w11092 = w11091 & w13597;
assign w11093 = (~w11092 & w9765) | (~w11092 & w13752) | (w9765 & w13752);
assign w11094 = ~w702 & ~w9783;
assign w11095 = ~w9780 & w11094;
assign w11096 = w9785 & ~w11095;
assign w11097 = (w9783 & w9780) | (w9783 & w13753) | (w9780 & w13753);
assign w11098 = ~w11096 & ~w11097;
assign w11099 = ~w688 & ~w9769;
assign w11100 = ~w9766 & w11099;
assign w11101 = w9771 & ~w11100;
assign w11102 = (w9769 & w9766) | (w9769 & w13754) | (w9766 & w13754);
assign w11103 = ~w11101 & ~w11102;
assign w11104 = ~w11098 & w11103;
assign w11105 = w11098 & ~w11103;
assign w11106 = ~w11104 & ~w11105;
assign w11107 = ~w11093 & ~w11106;
assign w11108 = ~w11092 & ~w11104;
assign w11109 = ~w11105 & w11108;
assign w11110 = ~w11090 & w11109;
assign w11111 = ~w11107 & ~w11110;
assign w11112 = ~w9743 & ~w9757;
assign w11113 = (~w11112 & w9728) | (~w11112 & w13598) | (w9728 & w13598);
assign w11114 = ~w9742 & ~w9756;
assign w11115 = w11114 & w13599;
assign w11116 = ~w11115 & ~w11113;
assign w11117 = ~w732 & ~w9747;
assign w11118 = ~w9744 & w11117;
assign w11119 = w9749 & ~w11118;
assign w11120 = (w9747 & w9744) | (w9747 & w13755) | (w9744 & w13755);
assign w11121 = ~w11119 & ~w11120;
assign w11122 = ~w757 & ~w9733;
assign w11123 = ~w9730 & w11122;
assign w11124 = w9735 & ~w11123;
assign w11125 = (w9733 & w9730) | (w9733 & w13756) | (w9730 & w13756);
assign w11126 = ~w11124 & ~w11125;
assign w11127 = ~w11121 & w11126;
assign w11128 = w11121 & ~w11126;
assign w11129 = ~w11127 & ~w11128;
assign w11130 = ~w11116 & ~w11129;
assign w11131 = ~w11115 & ~w11127;
assign w11132 = ~w11128 & w11131;
assign w11133 = ~w11113 & w11132;
assign w11134 = ~w11130 & ~w11133;
assign w11135 = ~w11111 & w11134;
assign w11136 = w11111 & ~w11134;
assign w11137 = ~w11135 & ~w11136;
assign w11138 = ~w11088 & ~w11137;
assign w11139 = w11088 & w11137;
assign w11140 = ~w11138 & ~w11139;
assign w11141 = ~w11084 & w11140;
assign w11142 = w11084 & ~w11140;
assign w11143 = ~w11141 & ~w11142;
assign w11144 = ~w11028 & ~w11143;
assign w11145 = w11028 & w11143;
assign w11146 = ~w11144 & ~w11145;
assign w11147 = ~w11024 & w11146;
assign w11148 = w11024 & ~w11146;
assign w11149 = ~w11147 & ~w11148;
assign w11150 = ~w10902 & ~w11149;
assign w11151 = w10902 & w11149;
assign w11152 = ~w11150 & ~w11151;
assign w11153 = ~w9547 & ~w9715;
assign w11154 = ~w9379 & ~w11153;
assign w11155 = w9547 & w9715;
assign w11156 = ~w11154 & ~w11155;
assign w11157 = ~w9629 & ~w9709;
assign w11158 = ~w9549 & ~w11157;
assign w11159 = w9629 & w9709;
assign w11160 = ~w11158 & ~w11159;
assign w11161 = ~w9667 & ~w9703;
assign w11162 = ~w9631 & ~w11161;
assign w11163 = w9667 & w9703;
assign w11164 = ~w11162 & ~w11163;
assign w11165 = ~w9683 & ~w9697;
assign w11166 = ~w9669 & ~w11165;
assign w11167 = ~w9682 & ~w9696;
assign w11168 = w11167 & w13600;
assign w11169 = (~w11168 & w9669) | (~w11168 & w13757) | (w9669 & w13757);
assign w11170 = ~w2900 & ~w9687;
assign w11171 = ~w9684 & w11170;
assign w11172 = w9689 & ~w11171;
assign w11173 = (w9687 & w9684) | (w9687 & w13758) | (w9684 & w13758);
assign w11174 = ~w11172 & ~w11173;
assign w11175 = ~w2886 & ~w9673;
assign w11176 = ~w9670 & w11175;
assign w11177 = w9675 & ~w11176;
assign w11178 = (w9673 & w9670) | (w9673 & w13759) | (w9670 & w13759);
assign w11179 = ~w11177 & ~w11178;
assign w11180 = ~w11174 & w11179;
assign w11181 = w11174 & ~w11179;
assign w11182 = ~w11180 & ~w11181;
assign w11183 = ~w11169 & ~w11182;
assign w11184 = ~w11168 & ~w11180;
assign w11185 = ~w11181 & w11184;
assign w11186 = ~w11166 & w11185;
assign w11187 = ~w11183 & ~w11186;
assign w11188 = ~w9647 & ~w9661;
assign w11189 = (~w11188 & w9632) | (~w11188 & w13601) | (w9632 & w13601);
assign w11190 = ~w9646 & ~w9660;
assign w11191 = w11190 & w13602;
assign w11192 = ~w11191 & ~w11189;
assign w11193 = ~w2838 & ~w9651;
assign w11194 = ~w9648 & w11193;
assign w11195 = w9653 & ~w11194;
assign w11196 = (w9651 & w9648) | (w9651 & w13760) | (w9648 & w13760);
assign w11197 = ~w11195 & ~w11196;
assign w11198 = ~w2863 & ~w9637;
assign w11199 = ~w9634 & w11198;
assign w11200 = w9639 & ~w11199;
assign w11201 = (w9637 & w9634) | (w9637 & w13761) | (w9634 & w13761);
assign w11202 = ~w11200 & ~w11201;
assign w11203 = ~w11197 & w11202;
assign w11204 = w11197 & ~w11202;
assign w11205 = ~w11203 & ~w11204;
assign w11206 = ~w11192 & ~w11205;
assign w11207 = ~w11191 & ~w11203;
assign w11208 = ~w11204 & w11207;
assign w11209 = ~w11189 & w11208;
assign w11210 = ~w11206 & ~w11209;
assign w11211 = ~w11187 & w11210;
assign w11212 = w11187 & ~w11210;
assign w11213 = ~w11211 & ~w11212;
assign w11214 = ~w11164 & ~w11213;
assign w11215 = w11164 & w11213;
assign w11216 = ~w11214 & ~w11215;
assign w11217 = ~w9587 & ~w9623;
assign w11218 = ~w9551 & ~w11217;
assign w11219 = w9587 & w9623;
assign w11220 = ~w11218 & ~w11219;
assign w11221 = ~w9603 & ~w9617;
assign w11222 = ~w9589 & ~w11221;
assign w11223 = ~w9602 & ~w9616;
assign w11224 = w11223 & w13603;
assign w11225 = (~w11224 & w9589) | (~w11224 & w13762) | (w9589 & w13762);
assign w11226 = ~w2758 & ~w9607;
assign w11227 = ~w9604 & w11226;
assign w11228 = w9609 & ~w11227;
assign w11229 = (w9607 & w9604) | (w9607 & w13763) | (w9604 & w13763);
assign w11230 = ~w11228 & ~w11229;
assign w11231 = ~w2744 & ~w9593;
assign w11232 = ~w9590 & w11231;
assign w11233 = w9595 & ~w11232;
assign w11234 = (w9593 & w9590) | (w9593 & w13764) | (w9590 & w13764);
assign w11235 = ~w11233 & ~w11234;
assign w11236 = ~w11230 & w11235;
assign w11237 = w11230 & ~w11235;
assign w11238 = ~w11236 & ~w11237;
assign w11239 = ~w11225 & ~w11238;
assign w11240 = ~w11224 & ~w11236;
assign w11241 = ~w11237 & w11240;
assign w11242 = ~w11222 & w11241;
assign w11243 = ~w11239 & ~w11242;
assign w11244 = ~w9567 & ~w9581;
assign w11245 = (~w11244 & w9552) | (~w11244 & w13604) | (w9552 & w13604);
assign w11246 = ~w9566 & ~w9580;
assign w11247 = w11246 & w13605;
assign w11248 = ~w11247 & ~w11245;
assign w11249 = ~w2788 & ~w9571;
assign w11250 = ~w9568 & w11249;
assign w11251 = w9573 & ~w11250;
assign w11252 = (w9571 & w9568) | (w9571 & w13765) | (w9568 & w13765);
assign w11253 = ~w11251 & ~w11252;
assign w11254 = ~w2813 & ~w9557;
assign w11255 = ~w9554 & w11254;
assign w11256 = w9559 & ~w11255;
assign w11257 = (w9557 & w9554) | (w9557 & w13766) | (w9554 & w13766);
assign w11258 = ~w11256 & ~w11257;
assign w11259 = ~w11253 & w11258;
assign w11260 = w11253 & ~w11258;
assign w11261 = ~w11259 & ~w11260;
assign w11262 = ~w11248 & ~w11261;
assign w11263 = ~w11247 & ~w11259;
assign w11264 = ~w11260 & w11263;
assign w11265 = ~w11245 & w11264;
assign w11266 = ~w11262 & ~w11265;
assign w11267 = ~w11243 & w11266;
assign w11268 = w11243 & ~w11266;
assign w11269 = ~w11267 & ~w11268;
assign w11270 = ~w11220 & ~w11269;
assign w11271 = w11220 & w11269;
assign w11272 = ~w11270 & ~w11271;
assign w11273 = ~w11216 & w11272;
assign w11274 = w11216 & ~w11272;
assign w11275 = ~w11273 & ~w11274;
assign w11276 = ~w11160 & ~w11275;
assign w11277 = w11160 & w11275;
assign w11278 = ~w11276 & ~w11277;
assign w11279 = ~w9461 & ~w9541;
assign w11280 = ~w9381 & ~w11279;
assign w11281 = w9461 & w9541;
assign w11282 = ~w11280 & ~w11281;
assign w11283 = ~w9499 & ~w9535;
assign w11284 = ~w9463 & ~w11283;
assign w11285 = w9499 & w9535;
assign w11286 = ~w11284 & ~w11285;
assign w11287 = ~w9515 & ~w9529;
assign w11288 = ~w9501 & ~w11287;
assign w11289 = ~w9514 & ~w9528;
assign w11290 = w11289 & w13606;
assign w11291 = (~w11290 & w9501) | (~w11290 & w13767) | (w9501 & w13767);
assign w11292 = ~w3015 & ~w9519;
assign w11293 = ~w9516 & w11292;
assign w11294 = w9521 & ~w11293;
assign w11295 = (w9519 & w9516) | (w9519 & w13768) | (w9516 & w13768);
assign w11296 = ~w11294 & ~w11295;
assign w11297 = ~w3001 & ~w9505;
assign w11298 = ~w9502 & w11297;
assign w11299 = w9507 & ~w11298;
assign w11300 = (w9505 & w9502) | (w9505 & w13769) | (w9502 & w13769);
assign w11301 = ~w11299 & ~w11300;
assign w11302 = ~w11296 & w11301;
assign w11303 = w11296 & ~w11301;
assign w11304 = ~w11302 & ~w11303;
assign w11305 = ~w11291 & ~w11304;
assign w11306 = ~w11290 & ~w11302;
assign w11307 = ~w11303 & w11306;
assign w11308 = ~w11288 & w11307;
assign w11309 = ~w11305 & ~w11308;
assign w11310 = ~w9479 & ~w9493;
assign w11311 = (~w11310 & w9464) | (~w11310 & w13607) | (w9464 & w13607);
assign w11312 = ~w9478 & ~w9492;
assign w11313 = w11312 & w13608;
assign w11314 = ~w11313 & ~w11311;
assign w11315 = ~w2953 & ~w9483;
assign w11316 = ~w9480 & w11315;
assign w11317 = w9485 & ~w11316;
assign w11318 = (w9483 & w9480) | (w9483 & w13770) | (w9480 & w13770);
assign w11319 = ~w11317 & ~w11318;
assign w11320 = ~w2978 & ~w9469;
assign w11321 = ~w9466 & w11320;
assign w11322 = w9471 & ~w11321;
assign w11323 = (w9469 & w9466) | (w9469 & w13771) | (w9466 & w13771);
assign w11324 = ~w11322 & ~w11323;
assign w11325 = ~w11319 & w11324;
assign w11326 = w11319 & ~w11324;
assign w11327 = ~w11325 & ~w11326;
assign w11328 = ~w11314 & ~w11327;
assign w11329 = ~w11313 & ~w11325;
assign w11330 = ~w11326 & w11329;
assign w11331 = ~w11311 & w11330;
assign w11332 = ~w11328 & ~w11331;
assign w11333 = ~w11309 & w11332;
assign w11334 = w11309 & ~w11332;
assign w11335 = ~w11333 & ~w11334;
assign w11336 = ~w11286 & ~w11335;
assign w11337 = w11286 & w11335;
assign w11338 = ~w11336 & ~w11337;
assign w11339 = ~w9419 & ~w9455;
assign w11340 = ~w9383 & ~w11339;
assign w11341 = w9419 & w9455;
assign w11342 = ~w11340 & ~w11341;
assign w11343 = ~w9435 & ~w9449;
assign w11344 = ~w9421 & ~w11343;
assign w11345 = ~w9434 & ~w9448;
assign w11346 = w11345 & w13609;
assign w11347 = (~w11346 & w9421) | (~w11346 & w13772) | (w9421 & w13772);
assign w11348 = ~w3074 & ~w9439;
assign w11349 = ~w9436 & w11348;
assign w11350 = w9441 & ~w11349;
assign w11351 = (w9439 & w9436) | (w9439 & w13773) | (w9436 & w13773);
assign w11352 = ~w11350 & ~w11351;
assign w11353 = ~w3060 & ~w9425;
assign w11354 = ~w9422 & w11353;
assign w11355 = w9427 & ~w11354;
assign w11356 = (w9425 & w9422) | (w9425 & w13774) | (w9422 & w13774);
assign w11357 = ~w11355 & ~w11356;
assign w11358 = ~w11352 & w11357;
assign w11359 = w11352 & ~w11357;
assign w11360 = ~w11358 & ~w11359;
assign w11361 = ~w11347 & ~w11360;
assign w11362 = ~w11346 & ~w11358;
assign w11363 = ~w11359 & w11362;
assign w11364 = ~w11344 & w11363;
assign w11365 = ~w11361 & ~w11364;
assign w11366 = ~w9399 & ~w9413;
assign w11367 = (~w11366 & w9384) | (~w11366 & w13610) | (w9384 & w13610);
assign w11368 = ~w9398 & ~w9412;
assign w11369 = w11368 & w13611;
assign w11370 = ~w11369 & ~w11367;
assign w11371 = ~w3104 & ~w9403;
assign w11372 = ~w9400 & w11371;
assign w11373 = w9405 & ~w11372;
assign w11374 = (w9403 & w9400) | (w9403 & w13775) | (w9400 & w13775);
assign w11375 = ~w11373 & ~w11374;
assign w11376 = ~w3129 & ~w9389;
assign w11377 = ~w9386 & w11376;
assign w11378 = w9391 & ~w11377;
assign w11379 = (w9389 & w9386) | (w9389 & w13776) | (w9386 & w13776);
assign w11380 = ~w11378 & ~w11379;
assign w11381 = ~w11375 & w11380;
assign w11382 = w11375 & ~w11380;
assign w11383 = ~w11381 & ~w11382;
assign w11384 = ~w11370 & ~w11383;
assign w11385 = ~w11369 & ~w11381;
assign w11386 = ~w11382 & w11385;
assign w11387 = ~w11367 & w11386;
assign w11388 = ~w11384 & ~w11387;
assign w11389 = ~w11365 & w11388;
assign w11390 = w11365 & ~w11388;
assign w11391 = ~w11389 & ~w11390;
assign w11392 = ~w11342 & ~w11391;
assign w11393 = w11342 & w11391;
assign w11394 = ~w11392 & ~w11393;
assign w11395 = ~w11338 & w11394;
assign w11396 = w11338 & ~w11394;
assign w11397 = ~w11395 & ~w11396;
assign w11398 = ~w11282 & ~w11397;
assign w11399 = w11282 & w11397;
assign w11400 = ~w11398 & ~w11399;
assign w11401 = ~w11278 & w11400;
assign w11402 = w11278 & ~w11400;
assign w11403 = ~w11401 & ~w11402;
assign w11404 = ~w11156 & ~w11403;
assign w11405 = w11156 & w11403;
assign w11406 = ~w11404 & ~w11405;
assign w11407 = ~w11152 & w11406;
assign w11408 = w11152 & ~w11406;
assign w11409 = ~w11407 & ~w11408;
assign w11410 = ~w10898 & ~w11409;
assign w11411 = w10898 & w11409;
assign w11412 = ~w11410 & ~w11411;
assign w11413 = ~w10894 & ~w11412;
assign w11414 = (w11412 & w10891) | (w11412 & w13914) | (w10891 & w13914);
assign w11415 = ~w10893 & w11414;
assign w11416 = (~w11415 & w10075) | (~w11415 & w13432) | (w10075 & w13432);
assign w11417 = ~w10585 & ~w10888;
assign w11418 = w10585 & w10888;
assign w11419 = (~w11418 & w10078) | (~w11418 & w13433) | (w10078 & w13433);
assign w11420 = ~w10760 & ~w10881;
assign w11421 = (w10881 & w10757) | (w10881 & w13915) | (w10757 & w13915);
assign w11422 = ~w10759 & w11421;
assign w11423 = (~w11422 & w10590) | (~w11422 & w13434) | (w10590 & w13434);
assign w11424 = ~w10699 & ~w10753;
assign w11425 = ~w10697 & w10753;
assign w11426 = ~w10698 & w11425;
assign w11427 = (~w11426 & w10594) | (~w11426 & w13435) | (w10594 & w13435);
assign w11428 = ~w10652 & ~w10693;
assign w11429 = w10652 & w10693;
assign w11430 = (~w11429 & w10597) | (~w11429 & w13436) | (w10597 & w13436);
assign w11431 = ~w10656 & ~w10688;
assign w11432 = (~w10689 & w10656) | (~w10689 & w13437) | (w10656 & w13437);
assign w11433 = w10674 & w10679;
assign w11434 = (~w11433 & w10667) | (~w11433 & w12952) | (w10667 & w12952);
assign w11435 = ~w10674 & ~w10679;
assign w11436 = (~w11435 & w10660) | (~w11435 & w13916) | (w10660 & w13916);
assign w11437 = ~w11434 & w11436;
assign w11438 = ~w11435 & ~w11434;
assign w11439 = w10662 & ~w11438;
assign w11440 = ~w11437 & ~w11439;
assign w11441 = ~w11432 & w11440;
assign w11442 = ~w10689 & ~w11440;
assign w11443 = ~w11431 & w11442;
assign w11444 = ~w11441 & ~w11443;
assign w11445 = ~w10623 & ~w10646;
assign w11446 = ~w10600 & ~w11445;
assign w11447 = ~w10622 & ~w10645;
assign w11448 = w11447 & w13120;
assign w11449 = (~w11448 & w10600) | (~w11448 & w13438) | (w10600 & w13438);
assign w11450 = w10610 & w10615;
assign w11451 = ~w10605 & ~w11450;
assign w11452 = ~w10610 & ~w10615;
assign w11453 = (~w11452 & w10605) | (~w11452 & w13439) | (w10605 & w13439);
assign w11454 = w10633 & w10638;
assign w11455 = ~w10633 & ~w10638;
assign w11456 = (~w11455 & w10628) | (~w11455 & w13440) | (w10628 & w13440);
assign w11457 = ~w11453 & w11456;
assign w11458 = w11453 & ~w11456;
assign w11459 = ~w11457 & ~w11458;
assign w11460 = ~w11449 & ~w11459;
assign w11461 = ~w11448 & w11459;
assign w11462 = ~w11446 & w11461;
assign w11463 = ~w11460 & ~w11462;
assign w11464 = ~w11444 & w11463;
assign w11465 = w11444 & ~w11463;
assign w11466 = ~w11464 & ~w11465;
assign w11467 = w11430 & w11466;
assign w11468 = ~w11430 & ~w11466;
assign w11469 = ~w10725 & ~w10747;
assign w11470 = ~w10703 & ~w11469;
assign w11471 = ~w10724 & ~w10746;
assign w11472 = w11471 & w13917;
assign w11473 = w10712 & w10717;
assign w11474 = (~w11473 & w10705) | (~w11473 & w13918) | (w10705 & w13918);
assign w11475 = ~w10712 & ~w10717;
assign w11476 = ~w11475 & ~w11474;
assign w11477 = w10734 & w10739;
assign w11478 = ~w10734 & ~w10739;
assign w11479 = ~w11478 & w14068;
assign w11480 = ~w11476 & w11479;
assign w11481 = w11476 & ~w11479;
assign w11482 = ~w11480 & ~w11481;
assign w11483 = (~w11482 & w11470) | (~w11482 & w13920) | (w11470 & w13920);
assign w11484 = ~w11472 & w11482;
assign w11485 = ~w11470 & w11484;
assign w11486 = ~w11483 & ~w11485;
assign w11487 = ~w11468 & ~w11486;
assign w11488 = ~w11467 & w11487;
assign w11489 = ~w11467 & ~w11468;
assign w11490 = w11486 & ~w11489;
assign w11491 = ~w11488 & ~w11490;
assign w11492 = w11427 & w11491;
assign w11493 = ~w11427 & ~w11491;
assign w11494 = ~w10820 & ~w10875;
assign w11495 = w10820 & w10875;
assign w11496 = (~w11495 & w10764) | (~w11495 & w13921) | (w10764 & w13921);
assign w11497 = ~w10846 & ~w10869;
assign w11498 = ~w10823 & ~w11497;
assign w11499 = ~w10845 & ~w10868;
assign w11500 = w11499 & w13922;
assign w11501 = w10833 & w10838;
assign w11502 = ~w10828 & ~w11501;
assign w11503 = ~w10833 & ~w10838;
assign w11504 = (~w11503 & w10828) | (~w11503 & w13923) | (w10828 & w13923);
assign w11505 = w10856 & w10861;
assign w11506 = ~w10856 & ~w10861;
assign w11507 = (~w11506 & w10851) | (~w11506 & w13924) | (w10851 & w13924);
assign w11508 = ~w11504 & w11507;
assign w11509 = w11504 & ~w11507;
assign w11510 = ~w11508 & ~w11509;
assign w11511 = (~w11510 & w11498) | (~w11510 & w13925) | (w11498 & w13925);
assign w11512 = ~w11500 & w11510;
assign w11513 = ~w11498 & w11512;
assign w11514 = ~w11511 & ~w11513;
assign w11515 = ~w10791 & ~w10814;
assign w11516 = ~w10768 & ~w11515;
assign w11517 = ~w10790 & ~w10813;
assign w11518 = w11517 & w13926;
assign w11519 = w10778 & w10783;
assign w11520 = ~w10773 & ~w11519;
assign w11521 = ~w10778 & ~w10783;
assign w11522 = (~w11521 & w10773) | (~w11521 & w13927) | (w10773 & w13927);
assign w11523 = w10801 & w10806;
assign w11524 = ~w10801 & ~w10806;
assign w11525 = (~w11524 & w10796) | (~w11524 & w13928) | (w10796 & w13928);
assign w11526 = ~w11522 & w11525;
assign w11527 = w11522 & ~w11525;
assign w11528 = ~w11526 & ~w11527;
assign w11529 = (~w11528 & w11516) | (~w11528 & w13929) | (w11516 & w13929);
assign w11530 = ~w11518 & w11528;
assign w11531 = ~w11516 & w11530;
assign w11532 = ~w11529 & ~w11531;
assign w11533 = ~w11514 & w11532;
assign w11534 = w11514 & ~w11532;
assign w11535 = ~w11533 & ~w11534;
assign w11536 = ~w11496 & ~w11535;
assign w11537 = w11496 & w11535;
assign w11538 = ~w11536 & ~w11537;
assign w11539 = ~w11493 & ~w11538;
assign w11540 = ~w11492 & w11539;
assign w11541 = ~w11492 & ~w11493;
assign w11542 = w11538 & ~w11541;
assign w11543 = ~w11540 & ~w11542;
assign w11544 = ~w11423 & ~w11543;
assign w11545 = w11423 & w11543;
assign w11546 = ~w11544 & ~w11545;
assign w11547 = ~w10332 & ~w10579;
assign w11548 = w10332 & w10579;
assign w11549 = (~w11548 & w10082) | (~w11548 & w13441) | (w10082 & w13441);
assign w11550 = ~w10454 & ~w10573;
assign w11551 = w10454 & w10573;
assign w11552 = (~w11551 & w10335) | (~w11551 & w13442) | (w10335 & w13442);
assign w11553 = ~w10512 & ~w10567;
assign w11554 = w10512 & w10567;
assign w11555 = (~w11554 & w10457) | (~w11554 & w13443) | (w10457 & w13443);
assign w11556 = ~w10538 & ~w10561;
assign w11557 = ~w10515 & ~w11556;
assign w11558 = ~w10537 & ~w10560;
assign w11559 = w11558 & w13121;
assign w11560 = (~w11559 & w10515) | (~w11559 & w13444) | (w10515 & w13444);
assign w11561 = w10525 & w10530;
assign w11562 = ~w10520 & ~w11561;
assign w11563 = ~w10525 & ~w10530;
assign w11564 = (~w11563 & w10520) | (~w11563 & w13445) | (w10520 & w13445);
assign w11565 = w10548 & w10553;
assign w11566 = ~w10548 & ~w10553;
assign w11567 = (~w11566 & w10543) | (~w11566 & w13446) | (w10543 & w13446);
assign w11568 = ~w11564 & w11567;
assign w11569 = w11564 & ~w11567;
assign w11570 = ~w11568 & ~w11569;
assign w11571 = ~w11560 & ~w11570;
assign w11572 = ~w11559 & w11570;
assign w11573 = ~w11557 & w11572;
assign w11574 = ~w11571 & ~w11573;
assign w11575 = ~w10483 & ~w10506;
assign w11576 = ~w10460 & ~w11575;
assign w11577 = ~w10482 & ~w10505;
assign w11578 = w11577 & w13122;
assign w11579 = (~w11578 & w10460) | (~w11578 & w13447) | (w10460 & w13447);
assign w11580 = w10470 & w10475;
assign w11581 = ~w10465 & ~w11580;
assign w11582 = ~w10470 & ~w10475;
assign w11583 = (~w11582 & w10465) | (~w11582 & w13448) | (w10465 & w13448);
assign w11584 = w10493 & w10498;
assign w11585 = ~w10493 & ~w10498;
assign w11586 = (~w11585 & w10488) | (~w11585 & w13449) | (w10488 & w13449);
assign w11587 = ~w11583 & w11586;
assign w11588 = w11583 & ~w11586;
assign w11589 = ~w11587 & ~w11588;
assign w11590 = ~w11579 & ~w11589;
assign w11591 = ~w11578 & w11589;
assign w11592 = ~w11576 & w11591;
assign w11593 = ~w11590 & ~w11592;
assign w11594 = ~w11574 & w11593;
assign w11595 = w11574 & ~w11593;
assign w11596 = ~w11594 & ~w11595;
assign w11597 = ~w11555 & ~w11596;
assign w11598 = w11555 & w11596;
assign w11599 = ~w11597 & ~w11598;
assign w11600 = ~w10393 & ~w10448;
assign w11601 = w10393 & w10448;
assign w11602 = (~w11601 & w10338) | (~w11601 & w13450) | (w10338 & w13450);
assign w11603 = ~w10419 & ~w10442;
assign w11604 = ~w10396 & ~w11603;
assign w11605 = ~w10418 & ~w10441;
assign w11606 = w11605 & w13123;
assign w11607 = (~w11606 & w10396) | (~w11606 & w13451) | (w10396 & w13451);
assign w11608 = w10406 & w10411;
assign w11609 = ~w10401 & ~w11608;
assign w11610 = ~w10406 & ~w10411;
assign w11611 = (~w11610 & w10401) | (~w11610 & w13452) | (w10401 & w13452);
assign w11612 = w10429 & w10434;
assign w11613 = ~w10429 & ~w10434;
assign w11614 = (~w11613 & w10424) | (~w11613 & w13453) | (w10424 & w13453);
assign w11615 = ~w11611 & w11614;
assign w11616 = w11611 & ~w11614;
assign w11617 = ~w11615 & ~w11616;
assign w11618 = ~w11607 & ~w11617;
assign w11619 = ~w11606 & w11617;
assign w11620 = ~w11604 & w11619;
assign w11621 = ~w11618 & ~w11620;
assign w11622 = ~w10364 & ~w10387;
assign w11623 = ~w10341 & ~w11622;
assign w11624 = ~w10363 & ~w10386;
assign w11625 = w11624 & w13124;
assign w11626 = (~w11625 & w10341) | (~w11625 & w13454) | (w10341 & w13454);
assign w11627 = w10351 & w10356;
assign w11628 = ~w10346 & ~w11627;
assign w11629 = ~w10351 & ~w10356;
assign w11630 = (~w11629 & w10346) | (~w11629 & w13455) | (w10346 & w13455);
assign w11631 = w10374 & w10379;
assign w11632 = ~w10374 & ~w10379;
assign w11633 = (~w11632 & w10369) | (~w11632 & w13456) | (w10369 & w13456);
assign w11634 = ~w11630 & w11633;
assign w11635 = w11630 & ~w11633;
assign w11636 = ~w11634 & ~w11635;
assign w11637 = ~w11626 & ~w11636;
assign w11638 = ~w11625 & w11636;
assign w11639 = ~w11623 & w11638;
assign w11640 = ~w11637 & ~w11639;
assign w11641 = ~w11621 & w11640;
assign w11642 = w11621 & ~w11640;
assign w11643 = ~w11641 & ~w11642;
assign w11644 = ~w11602 & ~w11643;
assign w11645 = w11602 & w11643;
assign w11646 = ~w11644 & ~w11645;
assign w11647 = ~w11599 & w11646;
assign w11648 = w11599 & ~w11646;
assign w11649 = ~w11647 & ~w11648;
assign w11650 = ~w11552 & ~w11649;
assign w11651 = w11552 & w11649;
assign w11652 = ~w11650 & ~w11651;
assign w11653 = ~w10207 & ~w10326;
assign w11654 = w10207 & w10326;
assign w11655 = (~w11654 & w10086) | (~w11654 & w13457) | (w10086 & w13457);
assign w11656 = ~w10265 & ~w10320;
assign w11657 = w10265 & w10320;
assign w11658 = (~w11657 & w10210) | (~w11657 & w13458) | (w10210 & w13458);
assign w11659 = ~w10291 & ~w10314;
assign w11660 = ~w10268 & ~w11659;
assign w11661 = ~w10290 & ~w10313;
assign w11662 = w11661 & w13125;
assign w11663 = (~w11662 & w10268) | (~w11662 & w13459) | (w10268 & w13459);
assign w11664 = w10278 & w10283;
assign w11665 = ~w10273 & ~w11664;
assign w11666 = ~w10278 & ~w10283;
assign w11667 = (~w11666 & w10273) | (~w11666 & w13460) | (w10273 & w13460);
assign w11668 = w10301 & w10306;
assign w11669 = ~w10301 & ~w10306;
assign w11670 = (~w11669 & w10296) | (~w11669 & w13461) | (w10296 & w13461);
assign w11671 = ~w11667 & w11670;
assign w11672 = w11667 & ~w11670;
assign w11673 = ~w11671 & ~w11672;
assign w11674 = ~w11663 & ~w11673;
assign w11675 = ~w11662 & w11673;
assign w11676 = ~w11660 & w11675;
assign w11677 = ~w11674 & ~w11676;
assign w11678 = ~w10236 & ~w10259;
assign w11679 = ~w10213 & ~w11678;
assign w11680 = ~w10235 & ~w10258;
assign w11681 = w11680 & w13126;
assign w11682 = (~w11681 & w10213) | (~w11681 & w13462) | (w10213 & w13462);
assign w11683 = w10223 & w10228;
assign w11684 = ~w10218 & ~w11683;
assign w11685 = ~w10223 & ~w10228;
assign w11686 = (~w11685 & w10218) | (~w11685 & w13463) | (w10218 & w13463);
assign w11687 = w10246 & w10251;
assign w11688 = ~w10246 & ~w10251;
assign w11689 = (~w11688 & w10241) | (~w11688 & w13464) | (w10241 & w13464);
assign w11690 = ~w11686 & w11689;
assign w11691 = w11686 & ~w11689;
assign w11692 = ~w11690 & ~w11691;
assign w11693 = ~w11682 & ~w11692;
assign w11694 = ~w11681 & w11692;
assign w11695 = ~w11679 & w11694;
assign w11696 = ~w11693 & ~w11695;
assign w11697 = ~w11677 & w11696;
assign w11698 = w11677 & ~w11696;
assign w11699 = ~w11697 & ~w11698;
assign w11700 = ~w11658 & ~w11699;
assign w11701 = w11658 & w11699;
assign w11702 = ~w11700 & ~w11701;
assign w11703 = ~w10146 & ~w10201;
assign w11704 = w10146 & w10201;
assign w11705 = (~w11704 & w10090) | (~w11704 & w13465) | (w10090 & w13465);
assign w11706 = ~w10172 & ~w10195;
assign w11707 = ~w10149 & ~w11706;
assign w11708 = ~w10171 & ~w10194;
assign w11709 = w11708 & w13127;
assign w11710 = (~w11709 & w10149) | (~w11709 & w13466) | (w10149 & w13466);
assign w11711 = w10159 & w10164;
assign w11712 = ~w10154 & ~w11711;
assign w11713 = ~w10159 & ~w10164;
assign w11714 = (~w11713 & w10154) | (~w11713 & w13467) | (w10154 & w13467);
assign w11715 = w10182 & w10187;
assign w11716 = ~w10182 & ~w10187;
assign w11717 = (~w11716 & w10177) | (~w11716 & w13468) | (w10177 & w13468);
assign w11718 = ~w11714 & w11717;
assign w11719 = w11714 & ~w11717;
assign w11720 = ~w11718 & ~w11719;
assign w11721 = ~w11710 & ~w11720;
assign w11722 = ~w11709 & w11720;
assign w11723 = ~w11707 & w11722;
assign w11724 = ~w11721 & ~w11723;
assign w11725 = ~w10117 & ~w10140;
assign w11726 = ~w10094 & ~w11725;
assign w11727 = ~w10116 & ~w10139;
assign w11728 = w11727 & w13128;
assign w11729 = w10104 & w10109;
assign w11730 = ~w10099 & ~w11729;
assign w11731 = ~w10104 & ~w10109;
assign w11732 = (~w11731 & w10099) | (~w11731 & w13129) | (w10099 & w13129);
assign w11733 = w10127 & w10132;
assign w11734 = ~w10127 & ~w10132;
assign w11735 = (~w11734 & w10122) | (~w11734 & w13130) | (w10122 & w13130);
assign w11736 = ~w11732 & w11735;
assign w11737 = w11732 & ~w11735;
assign w11738 = ~w11736 & ~w11737;
assign w11739 = (~w11738 & w11726) | (~w11738 & w13131) | (w11726 & w13131);
assign w11740 = ~w11728 & w11738;
assign w11741 = ~w11726 & w11740;
assign w11742 = ~w11739 & ~w11741;
assign w11743 = ~w11724 & w11742;
assign w11744 = w11724 & ~w11742;
assign w11745 = ~w11743 & ~w11744;
assign w11746 = ~w11705 & ~w11745;
assign w11747 = w11705 & w11745;
assign w11748 = ~w11746 & ~w11747;
assign w11749 = ~w11702 & w11748;
assign w11750 = w11702 & ~w11748;
assign w11751 = ~w11749 & ~w11750;
assign w11752 = ~w11655 & ~w11751;
assign w11753 = w11655 & w11751;
assign w11754 = ~w11752 & ~w11753;
assign w11755 = ~w11652 & w11754;
assign w11756 = w11652 & ~w11754;
assign w11757 = ~w11755 & ~w11756;
assign w11758 = ~w11549 & ~w11757;
assign w11759 = w11549 & w11757;
assign w11760 = ~w11758 & ~w11759;
assign w11761 = ~w11546 & w11760;
assign w11762 = w11546 & ~w11760;
assign w11763 = ~w11761 & ~w11762;
assign w11764 = ~w11419 & ~w11763;
assign w11765 = w11419 & w11763;
assign w11766 = ~w11764 & ~w11765;
assign w11767 = ~w11152 & ~w11406;
assign w11768 = w11152 & w11406;
assign w11769 = (~w11768 & w10898) | (~w11768 & w13132) | (w10898 & w13132);
assign w11770 = ~w11278 & ~w11400;
assign w11771 = w11278 & w11400;
assign w11772 = (~w11771 & w11156) | (~w11771 & w13133) | (w11156 & w13133);
assign w11773 = ~w11338 & ~w11394;
assign w11774 = w11338 & w11394;
assign w11775 = (~w11774 & w11282) | (~w11774 & w13134) | (w11282 & w13134);
assign w11776 = ~w11365 & ~w11388;
assign w11777 = ~w11342 & ~w11776;
assign w11778 = ~w11364 & ~w11387;
assign w11779 = w11778 & w13777;
assign w11780 = (~w11779 & w11342) | (~w11779 & w13135) | (w11342 & w13135);
assign w11781 = w11352 & w11357;
assign w11782 = ~w11347 & ~w11781;
assign w11783 = ~w11352 & ~w11357;
assign w11784 = (~w11783 & w11347) | (~w11783 & w13930) | (w11347 & w13930);
assign w11785 = w11375 & w11380;
assign w11786 = ~w11375 & ~w11380;
assign w11787 = (~w11786 & w11370) | (~w11786 & w13931) | (w11370 & w13931);
assign w11788 = ~w11784 & w11787;
assign w11789 = w11784 & ~w11787;
assign w11790 = ~w11788 & ~w11789;
assign w11791 = ~w11780 & ~w11790;
assign w11792 = ~w11779 & w11790;
assign w11793 = ~w11777 & w11792;
assign w11794 = ~w11791 & ~w11793;
assign w11795 = ~w11309 & ~w11332;
assign w11796 = ~w11286 & ~w11795;
assign w11797 = ~w11308 & ~w11331;
assign w11798 = w11797 & w13778;
assign w11799 = (~w11798 & w11286) | (~w11798 & w13136) | (w11286 & w13136);
assign w11800 = w11296 & w11301;
assign w11801 = ~w11291 & ~w11800;
assign w11802 = ~w11296 & ~w11301;
assign w11803 = (~w11802 & w11291) | (~w11802 & w13932) | (w11291 & w13932);
assign w11804 = w11319 & w11324;
assign w11805 = ~w11319 & ~w11324;
assign w11806 = (~w11805 & w11314) | (~w11805 & w13933) | (w11314 & w13933);
assign w11807 = ~w11803 & w11806;
assign w11808 = w11803 & ~w11806;
assign w11809 = ~w11807 & ~w11808;
assign w11810 = ~w11799 & ~w11809;
assign w11811 = ~w11798 & w11809;
assign w11812 = ~w11796 & w11811;
assign w11813 = ~w11810 & ~w11812;
assign w11814 = ~w11794 & w11813;
assign w11815 = w11794 & ~w11813;
assign w11816 = ~w11814 & ~w11815;
assign w11817 = ~w11775 & ~w11816;
assign w11818 = w11775 & w11816;
assign w11819 = ~w11817 & ~w11818;
assign w11820 = ~w11216 & ~w11272;
assign w11821 = w11216 & w11272;
assign w11822 = (~w11821 & w11160) | (~w11821 & w13137) | (w11160 & w13137);
assign w11823 = ~w11243 & ~w11266;
assign w11824 = ~w11220 & ~w11823;
assign w11825 = ~w11242 & ~w11265;
assign w11826 = w11825 & w13779;
assign w11827 = (~w11826 & w11220) | (~w11826 & w13138) | (w11220 & w13138);
assign w11828 = w11230 & w11235;
assign w11829 = ~w11225 & ~w11828;
assign w11830 = ~w11230 & ~w11235;
assign w11831 = (~w11830 & w11225) | (~w11830 & w13934) | (w11225 & w13934);
assign w11832 = w11253 & w11258;
assign w11833 = ~w11253 & ~w11258;
assign w11834 = (~w11833 & w11248) | (~w11833 & w13935) | (w11248 & w13935);
assign w11835 = ~w11831 & w11834;
assign w11836 = w11831 & ~w11834;
assign w11837 = ~w11835 & ~w11836;
assign w11838 = ~w11827 & ~w11837;
assign w11839 = ~w11826 & w11837;
assign w11840 = ~w11824 & w11839;
assign w11841 = ~w11838 & ~w11840;
assign w11842 = ~w11187 & ~w11210;
assign w11843 = ~w11164 & ~w11842;
assign w11844 = ~w11186 & ~w11209;
assign w11845 = w11844 & w13780;
assign w11846 = (~w11845 & w11164) | (~w11845 & w13139) | (w11164 & w13139);
assign w11847 = w11174 & w11179;
assign w11848 = ~w11169 & ~w11847;
assign w11849 = ~w11174 & ~w11179;
assign w11850 = (~w11849 & w11169) | (~w11849 & w13936) | (w11169 & w13936);
assign w11851 = w11197 & w11202;
assign w11852 = ~w11197 & ~w11202;
assign w11853 = (~w11852 & w11192) | (~w11852 & w13937) | (w11192 & w13937);
assign w11854 = ~w11850 & w11853;
assign w11855 = w11850 & ~w11853;
assign w11856 = ~w11854 & ~w11855;
assign w11857 = ~w11846 & ~w11856;
assign w11858 = ~w11845 & w11856;
assign w11859 = ~w11843 & w11858;
assign w11860 = ~w11857 & ~w11859;
assign w11861 = ~w11841 & w11860;
assign w11862 = w11841 & ~w11860;
assign w11863 = ~w11861 & ~w11862;
assign w11864 = ~w11822 & ~w11863;
assign w11865 = w11822 & w11863;
assign w11866 = ~w11864 & ~w11865;
assign w11867 = ~w11819 & w11866;
assign w11868 = w11819 & ~w11866;
assign w11869 = ~w11867 & ~w11868;
assign w11870 = ~w11772 & ~w11869;
assign w11871 = w11772 & w11869;
assign w11872 = ~w11870 & ~w11871;
assign w11873 = ~w11024 & ~w11146;
assign w11874 = w11024 & w11146;
assign w11875 = (~w11874 & w10902) | (~w11874 & w13140) | (w10902 & w13140);
assign w11876 = ~w11084 & ~w11140;
assign w11877 = w11084 & w11140;
assign w11878 = (~w11877 & w11028) | (~w11877 & w13141) | (w11028 & w13141);
assign w11879 = ~w11111 & ~w11134;
assign w11880 = ~w11088 & ~w11879;
assign w11881 = ~w11110 & ~w11133;
assign w11882 = w11881 & w13781;
assign w11883 = (~w11882 & w11088) | (~w11882 & w13142) | (w11088 & w13142);
assign w11884 = w11098 & w11103;
assign w11885 = ~w11093 & ~w11884;
assign w11886 = ~w11098 & ~w11103;
assign w11887 = (~w11886 & w11093) | (~w11886 & w13938) | (w11093 & w13938);
assign w11888 = w11121 & w11126;
assign w11889 = ~w11121 & ~w11126;
assign w11890 = (~w11889 & w11116) | (~w11889 & w13939) | (w11116 & w13939);
assign w11891 = ~w11887 & w11890;
assign w11892 = w11887 & ~w11890;
assign w11893 = ~w11891 & ~w11892;
assign w11894 = ~w11883 & ~w11893;
assign w11895 = ~w11882 & w11893;
assign w11896 = ~w11880 & w11895;
assign w11897 = ~w11894 & ~w11896;
assign w11898 = ~w11055 & ~w11078;
assign w11899 = ~w11032 & ~w11898;
assign w11900 = ~w11054 & ~w11077;
assign w11901 = w11900 & w13782;
assign w11902 = (~w11901 & w11032) | (~w11901 & w13143) | (w11032 & w13143);
assign w11903 = w11042 & w11047;
assign w11904 = ~w11037 & ~w11903;
assign w11905 = ~w11042 & ~w11047;
assign w11906 = (~w11905 & w11037) | (~w11905 & w13940) | (w11037 & w13940);
assign w11907 = w11065 & w11070;
assign w11908 = ~w11065 & ~w11070;
assign w11909 = (~w11908 & w11060) | (~w11908 & w13941) | (w11060 & w13941);
assign w11910 = ~w11906 & w11909;
assign w11911 = w11906 & ~w11909;
assign w11912 = ~w11910 & ~w11911;
assign w11913 = ~w11902 & ~w11912;
assign w11914 = ~w11901 & w11912;
assign w11915 = ~w11899 & w11914;
assign w11916 = ~w11913 & ~w11915;
assign w11917 = ~w11897 & w11916;
assign w11918 = w11897 & ~w11916;
assign w11919 = ~w11917 & ~w11918;
assign w11920 = ~w11878 & ~w11919;
assign w11921 = w11878 & w11919;
assign w11922 = ~w11920 & ~w11921;
assign w11923 = ~w10962 & ~w11018;
assign w11924 = w10962 & w11018;
assign w11925 = (~w11924 & w10906) | (~w11924 & w13144) | (w10906 & w13144);
assign w11926 = ~w10989 & ~w11012;
assign w11927 = ~w10966 & ~w11926;
assign w11928 = ~w10988 & ~w11011;
assign w11929 = w11928 & w13783;
assign w11930 = (~w11929 & w10966) | (~w11929 & w13145) | (w10966 & w13145);
assign w11931 = w10976 & w10981;
assign w11932 = ~w10971 & ~w11931;
assign w11933 = ~w10976 & ~w10981;
assign w11934 = (~w11933 & w10971) | (~w11933 & w13942) | (w10971 & w13942);
assign w11935 = w10999 & w11004;
assign w11936 = ~w10999 & ~w11004;
assign w11937 = (~w11936 & w10994) | (~w11936 & w13943) | (w10994 & w13943);
assign w11938 = ~w11934 & w11937;
assign w11939 = w11934 & ~w11937;
assign w11940 = ~w11938 & ~w11939;
assign w11941 = ~w11930 & ~w11940;
assign w11942 = ~w11929 & w11940;
assign w11943 = ~w11927 & w11942;
assign w11944 = ~w11941 & ~w11943;
assign w11945 = ~w10933 & ~w10956;
assign w11946 = ~w10910 & ~w11945;
assign w11947 = ~w10932 & ~w10955;
assign w11948 = w11947 & w13784;
assign w11949 = (~w11948 & w10910) | (~w11948 & w13146) | (w10910 & w13146);
assign w11950 = w10920 & w10925;
assign w11951 = ~w10915 & ~w11950;
assign w11952 = ~w10920 & ~w10925;
assign w11953 = (~w11952 & w10915) | (~w11952 & w13944) | (w10915 & w13944);
assign w11954 = w10943 & w10948;
assign w11955 = ~w10943 & ~w10948;
assign w11956 = (~w11955 & w10938) | (~w11955 & w13945) | (w10938 & w13945);
assign w11957 = ~w11953 & w11956;
assign w11958 = w11953 & ~w11956;
assign w11959 = ~w11957 & ~w11958;
assign w11960 = ~w11949 & ~w11959;
assign w11961 = ~w11948 & w11959;
assign w11962 = ~w11946 & w11961;
assign w11963 = ~w11960 & ~w11962;
assign w11964 = ~w11944 & w11963;
assign w11965 = w11944 & ~w11963;
assign w11966 = ~w11964 & ~w11965;
assign w11967 = ~w11925 & ~w11966;
assign w11968 = w11925 & w11966;
assign w11969 = ~w11967 & ~w11968;
assign w11970 = ~w11922 & w11969;
assign w11971 = w11922 & ~w11969;
assign w11972 = ~w11970 & ~w11971;
assign w11973 = ~w11875 & ~w11972;
assign w11974 = w11875 & w11972;
assign w11975 = ~w11973 & ~w11974;
assign w11976 = ~w11872 & w11975;
assign w11977 = w11872 & ~w11975;
assign w11978 = ~w11976 & ~w11977;
assign w11979 = ~w11769 & ~w11978;
assign w11980 = w11769 & w11978;
assign w11981 = ~w11979 & ~w11980;
assign w11982 = ~w11766 & ~w11981;
assign w11983 = ~w11764 & w11981;
assign w11984 = ~w11765 & w11983;
assign w11985 = (~w11984 & w11416) | (~w11984 & w13147) | (w11416 & w13147);
assign w11986 = ~w11546 & ~w11760;
assign w11987 = w11546 & w11760;
assign w11988 = (~w11987 & w11419) | (~w11987 & w13148) | (w11419 & w13148);
assign w11989 = ~w11652 & ~w11754;
assign w11990 = w11652 & w11754;
assign w11991 = (~w11990 & w11549) | (~w11990 & w13149) | (w11549 & w13149);
assign w11992 = ~w11702 & ~w11748;
assign w11993 = w11702 & w11748;
assign w11994 = (~w11993 & w11655) | (~w11993 & w13150) | (w11655 & w13150);
assign w11995 = ~w11724 & ~w11742;
assign w11996 = ~w11705 & ~w11995;
assign w11997 = ~w11723 & ~w11741;
assign w11998 = w11997 & w13469;
assign w11999 = (~w11998 & w11705) | (~w11998 & w13151) | (w11705 & w13151);
assign w12000 = ~w11731 & ~w11734;
assign w12001 = (w12000 & w10122) | (w12000 & w13946) | (w10122 & w13946);
assign w12002 = ~w11730 & w12001;
assign w12003 = (~w12002 & w11726) | (~w12002 & w13152) | (w11726 & w13152);
assign w12004 = ~w11732 & ~w11735;
assign w12005 = (~w11726 & w13612) | (~w11726 & w13613) | (w13612 & w13613);
assign w12006 = ~w11713 & ~w11716;
assign w12007 = (w12006 & w10177) | (w12006 & w13947) | (w10177 & w13947);
assign w12008 = ~w11712 & w12007;
assign w12009 = ~w11714 & ~w11717;
assign w12010 = (~w11707 & w13614) | (~w11707 & w13615) | (w13614 & w13615);
assign w12011 = ~w12005 & w12010;
assign w12012 = w12005 & ~w12010;
assign w12013 = ~w12011 & ~w12012;
assign w12014 = ~w11999 & ~w12013;
assign w12015 = ~w11998 & w12013;
assign w12016 = ~w11996 & w12015;
assign w12017 = ~w12014 & ~w12016;
assign w12018 = ~w11677 & ~w11696;
assign w12019 = ~w11658 & ~w12018;
assign w12020 = ~w11676 & ~w11695;
assign w12021 = w12020 & w13470;
assign w12022 = (~w12021 & w11658) | (~w12021 & w13154) | (w11658 & w13154);
assign w12023 = ~w11685 & ~w11688;
assign w12024 = (w12023 & w10241) | (w12023 & w13948) | (w10241 & w13948);
assign w12025 = ~w11684 & w12024;
assign w12026 = (~w12025 & w11679) | (~w12025 & w13155) | (w11679 & w13155);
assign w12027 = ~w11686 & ~w11689;
assign w12028 = (~w11679 & w13616) | (~w11679 & w13617) | (w13616 & w13617);
assign w12029 = ~w11666 & ~w11669;
assign w12030 = (w12029 & w10296) | (w12029 & w13949) | (w10296 & w13949);
assign w12031 = ~w11665 & w12030;
assign w12032 = ~w11667 & ~w11670;
assign w12033 = (~w11660 & w13618) | (~w11660 & w13619) | (w13618 & w13619);
assign w12034 = ~w12028 & w12033;
assign w12035 = w12028 & ~w12033;
assign w12036 = ~w12034 & ~w12035;
assign w12037 = ~w12022 & ~w12036;
assign w12038 = ~w12021 & w12036;
assign w12039 = ~w12019 & w12038;
assign w12040 = ~w12037 & ~w12039;
assign w12041 = ~w12017 & w12040;
assign w12042 = w12017 & ~w12040;
assign w12043 = ~w12041 & ~w12042;
assign w12044 = ~w11994 & ~w12043;
assign w12045 = w11994 & w12043;
assign w12046 = ~w12044 & ~w12045;
assign w12047 = ~w11599 & ~w11646;
assign w12048 = w11599 & w11646;
assign w12049 = (~w12048 & w11552) | (~w12048 & w13157) | (w11552 & w13157);
assign w12050 = ~w11621 & ~w11640;
assign w12051 = ~w11602 & ~w12050;
assign w12052 = ~w11620 & ~w11639;
assign w12053 = w12052 & w13471;
assign w12054 = (~w12053 & w11602) | (~w12053 & w13158) | (w11602 & w13158);
assign w12055 = ~w11629 & ~w11632;
assign w12056 = (w12055 & w10369) | (w12055 & w13950) | (w10369 & w13950);
assign w12057 = ~w11628 & w12056;
assign w12058 = (~w12057 & w11623) | (~w12057 & w13159) | (w11623 & w13159);
assign w12059 = ~w11630 & ~w11633;
assign w12060 = (~w11623 & w13620) | (~w11623 & w13621) | (w13620 & w13621);
assign w12061 = ~w11610 & ~w11613;
assign w12062 = (w12061 & w10424) | (w12061 & w13951) | (w10424 & w13951);
assign w12063 = ~w11609 & w12062;
assign w12064 = ~w11611 & ~w11614;
assign w12065 = (~w11604 & w13622) | (~w11604 & w13623) | (w13622 & w13623);
assign w12066 = ~w12060 & w12065;
assign w12067 = w12060 & ~w12065;
assign w12068 = ~w12066 & ~w12067;
assign w12069 = ~w12054 & ~w12068;
assign w12070 = ~w12053 & w12068;
assign w12071 = ~w12051 & w12070;
assign w12072 = ~w12069 & ~w12071;
assign w12073 = ~w11574 & ~w11593;
assign w12074 = ~w11555 & ~w12073;
assign w12075 = ~w11573 & ~w11592;
assign w12076 = w12075 & w13472;
assign w12077 = (~w12076 & w11555) | (~w12076 & w13161) | (w11555 & w13161);
assign w12078 = ~w11582 & ~w11585;
assign w12079 = (w12078 & w10488) | (w12078 & w13952) | (w10488 & w13952);
assign w12080 = ~w11581 & w12079;
assign w12081 = (~w12080 & w11576) | (~w12080 & w13162) | (w11576 & w13162);
assign w12082 = ~w11583 & ~w11586;
assign w12083 = (~w11576 & w13624) | (~w11576 & w13625) | (w13624 & w13625);
assign w12084 = ~w11563 & ~w11566;
assign w12085 = (w12084 & w10543) | (w12084 & w13953) | (w10543 & w13953);
assign w12086 = ~w11562 & w12085;
assign w12087 = ~w11564 & ~w11567;
assign w12088 = (~w11557 & w13626) | (~w11557 & w13627) | (w13626 & w13627);
assign w12089 = ~w12083 & w12088;
assign w12090 = w12083 & ~w12088;
assign w12091 = ~w12089 & ~w12090;
assign w12092 = ~w12077 & ~w12091;
assign w12093 = ~w12076 & w12091;
assign w12094 = ~w12074 & w12093;
assign w12095 = ~w12092 & ~w12094;
assign w12096 = ~w12072 & w12095;
assign w12097 = w12072 & ~w12095;
assign w12098 = ~w12096 & ~w12097;
assign w12099 = ~w12049 & ~w12098;
assign w12100 = w12049 & w12098;
assign w12101 = ~w12099 & ~w12100;
assign w12102 = ~w12046 & w12101;
assign w12103 = w12046 & ~w12101;
assign w12104 = ~w12102 & ~w12103;
assign w12105 = ~w11991 & ~w12104;
assign w12106 = w11991 & w12104;
assign w12107 = ~w12105 & ~w12106;
assign w12108 = ~w11538 & ~w11541;
assign w12109 = ~w11493 & w11538;
assign w12110 = ~w11492 & w12109;
assign w12111 = (~w12110 & w11423) | (~w12110 & w13164) | (w11423 & w13164);
assign w12112 = ~w11486 & ~w11489;
assign w12113 = ~w11427 & ~w12112;
assign w12114 = ~w11468 & w11486;
assign w12115 = ~w11467 & w12114;
assign w12116 = (~w12115 & w11427) | (~w12115 & w13165) | (w11427 & w13165);
assign w12117 = ~w11444 & ~w11463;
assign w12118 = ~w11430 & ~w12117;
assign w12119 = ~w11443 & ~w11462;
assign w12120 = w12119 & w13473;
assign w12121 = (~w12120 & w11430) | (~w12120 & w13166) | (w11430 & w13166);
assign w12122 = ~w11452 & ~w11455;
assign w12123 = (w12122 & w10628) | (w12122 & w13785) | (w10628 & w13785);
assign w12124 = ~w11451 & w12123;
assign w12125 = (~w12124 & w11446) | (~w12124 & w13167) | (w11446 & w13167);
assign w12126 = ~w11453 & ~w11456;
assign w12127 = (~w11446 & w13628) | (~w11446 & w13629) | (w13628 & w13629);
assign w12128 = (~w11431 & w13630) | (~w11431 & w13631) | (w13630 & w13631);
assign w12129 = ~w12127 & w12128;
assign w12130 = w12127 & ~w12128;
assign w12131 = ~w12129 & ~w12130;
assign w12132 = ~w12121 & ~w12131;
assign w12133 = ~w12120 & w12131;
assign w12134 = ~w12118 & w12133;
assign w12135 = ~w11475 & ~w11478;
assign w12136 = w12135 & w14068;
assign w12137 = ~w11474 & w12136;
assign w12138 = ~w11476 & ~w11479;
assign w12139 = (~w11470 & w13954) | (~w11470 & w13955) | (w13954 & w13955);
assign w12140 = (w12139 & w12118) | (w12139 & w13632) | (w12118 & w13632);
assign w12141 = ~w12132 & w12140;
assign w12142 = ~w12132 & ~w12134;
assign w12143 = ~w12139 & ~w12142;
assign w12144 = ~w12141 & ~w12143;
assign w12145 = ~w12116 & ~w12144;
assign w12146 = ~w12115 & ~w12141;
assign w12147 = ~w12113 & w13633;
assign w12148 = ~w12145 & ~w12147;
assign w12149 = ~w11514 & ~w11532;
assign w12150 = ~w11496 & ~w12149;
assign w12151 = ~w11513 & ~w11531;
assign w12152 = w12151 & w13956;
assign w12153 = (~w12152 & w11496) | (~w12152 & w13169) | (w11496 & w13169);
assign w12154 = ~w11521 & ~w11524;
assign w12155 = (w12154 & w10796) | (w12154 & w13957) | (w10796 & w13957);
assign w12156 = ~w11520 & w12155;
assign w12157 = (~w12156 & w11516) | (~w12156 & w13958) | (w11516 & w13958);
assign w12158 = ~w11522 & ~w11525;
assign w12159 = (~w11516 & w13959) | (~w11516 & w13960) | (w13959 & w13960);
assign w12160 = ~w11503 & ~w11506;
assign w12161 = (w12160 & w10851) | (w12160 & w13961) | (w10851 & w13961);
assign w12162 = ~w11502 & w12161;
assign w12163 = ~w11504 & ~w11507;
assign w12164 = (~w11498 & w13963) | (~w11498 & w13964) | (w13963 & w13964);
assign w12165 = ~w12159 & w12164;
assign w12166 = w12159 & ~w12164;
assign w12167 = ~w12165 & ~w12166;
assign w12168 = ~w12153 & ~w12167;
assign w12169 = ~w12152 & w12167;
assign w12170 = ~w12150 & w12169;
assign w12171 = ~w12168 & ~w12170;
assign w12172 = (w12171 & w12147) | (w12171 & w13170) | (w12147 & w13170);
assign w12173 = ~w12145 & ~w12171;
assign w12174 = ~w12147 & w12173;
assign w12175 = ~w12172 & ~w12174;
assign w12176 = ~w12111 & ~w12175;
assign w12177 = w12111 & w12175;
assign w12178 = ~w12176 & ~w12177;
assign w12179 = ~w12107 & w12178;
assign w12180 = w12107 & ~w12178;
assign w12181 = ~w12179 & ~w12180;
assign w12182 = ~w11988 & ~w12181;
assign w12183 = w11988 & w12181;
assign w12184 = ~w12182 & ~w12183;
assign w12185 = ~w11872 & ~w11975;
assign w12186 = w11872 & w11975;
assign w12187 = (~w12186 & w11769) | (~w12186 & w13965) | (w11769 & w13965);
assign w12188 = ~w11922 & ~w11969;
assign w12189 = w11922 & w11969;
assign w12190 = (~w12189 & w11875) | (~w12189 & w13966) | (w11875 & w13966);
assign w12191 = ~w11944 & ~w11963;
assign w12192 = ~w11925 & ~w12191;
assign w12193 = ~w11943 & ~w11962;
assign w12194 = w12193 & w13967;
assign w12195 = ~w11952 & ~w11955;
assign w12196 = (w12195 & w10938) | (w12195 & w13968) | (w10938 & w13968);
assign w12197 = ~w11951 & w12196;
assign w12198 = ~w11949 & ~w12197;
assign w12199 = ~w11953 & ~w11956;
assign w12200 = (~w12199 & w11949) | (~w12199 & w13969) | (w11949 & w13969);
assign w12201 = ~w11933 & ~w11936;
assign w12202 = (w12201 & w10994) | (w12201 & w13970) | (w10994 & w13970);
assign w12203 = ~w11932 & w12202;
assign w12204 = ~w11934 & ~w11937;
assign w12205 = (~w12204 & w11930) | (~w12204 & w13971) | (w11930 & w13971);
assign w12206 = ~w12200 & w12205;
assign w12207 = w12200 & ~w12205;
assign w12208 = ~w12206 & ~w12207;
assign w12209 = (~w12208 & w12192) | (~w12208 & w13972) | (w12192 & w13972);
assign w12210 = ~w12194 & w12208;
assign w12211 = ~w12192 & w12210;
assign w12212 = ~w12209 & ~w12211;
assign w12213 = ~w11897 & ~w11916;
assign w12214 = ~w11878 & ~w12213;
assign w12215 = ~w11896 & ~w11915;
assign w12216 = w12215 & w13973;
assign w12217 = ~w11905 & ~w11908;
assign w12218 = (w12217 & w11060) | (w12217 & w13974) | (w11060 & w13974);
assign w12219 = ~w11904 & w12218;
assign w12220 = ~w11902 & ~w12219;
assign w12221 = ~w11906 & ~w11909;
assign w12222 = (~w12221 & w11902) | (~w12221 & w13975) | (w11902 & w13975);
assign w12223 = ~w11886 & ~w11889;
assign w12224 = (w12223 & w11116) | (w12223 & w13976) | (w11116 & w13976);
assign w12225 = ~w11885 & w12224;
assign w12226 = ~w11887 & ~w11890;
assign w12227 = (~w12226 & w11883) | (~w12226 & w13977) | (w11883 & w13977);
assign w12228 = ~w12222 & w12227;
assign w12229 = w12222 & ~w12227;
assign w12230 = ~w12228 & ~w12229;
assign w12231 = (~w12230 & w12214) | (~w12230 & w13978) | (w12214 & w13978);
assign w12232 = ~w12216 & w12230;
assign w12233 = ~w12214 & w12232;
assign w12234 = ~w12231 & ~w12233;
assign w12235 = ~w12212 & w12234;
assign w12236 = w12212 & ~w12234;
assign w12237 = ~w12235 & ~w12236;
assign w12238 = ~w12190 & ~w12237;
assign w12239 = w12190 & w12237;
assign w12240 = ~w12238 & ~w12239;
assign w12241 = ~w11819 & ~w11866;
assign w12242 = w11819 & w11866;
assign w12243 = (~w12242 & w11772) | (~w12242 & w13979) | (w11772 & w13979);
assign w12244 = ~w11841 & ~w11860;
assign w12245 = ~w11822 & ~w12244;
assign w12246 = ~w11840 & ~w11859;
assign w12247 = w12246 & w13980;
assign w12248 = ~w11849 & ~w11852;
assign w12249 = (w12248 & w11192) | (w12248 & w13981) | (w11192 & w13981);
assign w12250 = ~w11848 & w12249;
assign w12251 = ~w11846 & ~w12250;
assign w12252 = ~w11850 & ~w11853;
assign w12253 = (~w12252 & w11846) | (~w12252 & w13982) | (w11846 & w13982);
assign w12254 = ~w11830 & ~w11833;
assign w12255 = (w12254 & w11248) | (w12254 & w13983) | (w11248 & w13983);
assign w12256 = ~w11829 & w12255;
assign w12257 = ~w11831 & ~w11834;
assign w12258 = (~w12257 & w11827) | (~w12257 & w13984) | (w11827 & w13984);
assign w12259 = ~w12253 & w12258;
assign w12260 = w12253 & ~w12258;
assign w12261 = ~w12259 & ~w12260;
assign w12262 = (~w12261 & w12245) | (~w12261 & w13985) | (w12245 & w13985);
assign w12263 = ~w12247 & w12261;
assign w12264 = ~w12245 & w12263;
assign w12265 = ~w12262 & ~w12264;
assign w12266 = ~w11794 & ~w11813;
assign w12267 = ~w11775 & ~w12266;
assign w12268 = ~w11793 & ~w11812;
assign w12269 = w12268 & w13986;
assign w12270 = ~w11802 & ~w11805;
assign w12271 = (w12270 & w11314) | (w12270 & w13987) | (w11314 & w13987);
assign w12272 = ~w11801 & w12271;
assign w12273 = ~w11799 & ~w12272;
assign w12274 = ~w11803 & ~w11806;
assign w12275 = (~w12274 & w11799) | (~w12274 & w13988) | (w11799 & w13988);
assign w12276 = ~w11783 & ~w11786;
assign w12277 = (w12276 & w11370) | (w12276 & w13989) | (w11370 & w13989);
assign w12278 = ~w11782 & w12277;
assign w12279 = ~w11784 & ~w11787;
assign w12280 = (~w12279 & w11780) | (~w12279 & w13990) | (w11780 & w13990);
assign w12281 = ~w12275 & w12280;
assign w12282 = w12275 & ~w12280;
assign w12283 = ~w12281 & ~w12282;
assign w12284 = (~w12283 & w12267) | (~w12283 & w13991) | (w12267 & w13991);
assign w12285 = ~w12269 & w12283;
assign w12286 = ~w12267 & w12285;
assign w12287 = ~w12284 & ~w12286;
assign w12288 = ~w12265 & w12287;
assign w12289 = w12265 & ~w12287;
assign w12290 = ~w12288 & ~w12289;
assign w12291 = ~w12243 & ~w12290;
assign w12292 = w12243 & w12290;
assign w12293 = ~w12291 & ~w12292;
assign w12294 = ~w12240 & w12293;
assign w12295 = w12240 & ~w12293;
assign w12296 = ~w12294 & ~w12295;
assign w12297 = ~w12187 & ~w12296;
assign w12298 = w12187 & w12296;
assign w12299 = ~w12297 & ~w12298;
assign w12300 = ~w12184 & ~w12299;
assign w12301 = ~w12182 & w12299;
assign w12302 = ~w12183 & w12301;
assign w12303 = (~w12302 & w11985) | (~w12302 & w13634) | (w11985 & w13634);
assign w12304 = ~w12107 & ~w12178;
assign w12305 = w12107 & w12178;
assign w12306 = (~w12305 & w11988) | (~w12305 & w13635) | (w11988 & w13635);
assign w12307 = ~w12148 & ~w12171;
assign w12308 = ~w12145 & w12171;
assign w12309 = ~w12147 & w12308;
assign w12310 = (~w12309 & w12111) | (~w12309 & w13636) | (w12111 & w13636);
assign w12311 = ~w12158 & ~w12163;
assign w12312 = w12311 & w14069;
assign w12313 = ~w12157 & w12312;
assign w12314 = ~w12159 & ~w12164;
assign w12315 = (~w12314 & w12153) | (~w12314 & w13992) | (w12153 & w13992);
assign w12316 = w12139 & ~w12142;
assign w12317 = (~w12139 & w12118) | (~w12139 & w13786) | (w12118 & w13786);
assign w12318 = ~w12132 & w12317;
assign w12319 = (~w12318 & w12116) | (~w12318 & w13637) | (w12116 & w13637);
assign w12320 = ~w11439 & ~w12126;
assign w12321 = w12320 & w14070;
assign w12322 = ~w12125 & w12321;
assign w12323 = ~w12127 & ~w12128;
assign w12324 = (~w12323 & w12121) | (~w12323 & w13993) | (w12121 & w13993);
assign w12325 = ~w12319 & w12324;
assign w12326 = ~w12318 & ~w12324;
assign w12327 = (w12326 & w12116) | (w12326 & w13787) | (w12116 & w13787);
assign w12328 = (~w12315 & w12325) | (~w12315 & w13788) | (w12325 & w13788);
assign w12329 = w12315 & ~w12327;
assign w12330 = ~w12325 & w12329;
assign w12331 = ~w12328 & ~w12330;
assign w12332 = ~w12310 & w12331;
assign w12333 = w12310 & ~w12331;
assign w12334 = ~w12332 & ~w12333;
assign w12335 = ~w12046 & ~w12101;
assign w12336 = w12046 & w12101;
assign w12337 = (~w12336 & w11991) | (~w12336 & w13638) | (w11991 & w13638);
assign w12338 = ~w12072 & ~w12095;
assign w12339 = ~w12049 & ~w12338;
assign w12340 = ~w12071 & ~w12094;
assign w12341 = w12340 & w13171;
assign w12342 = (~w12341 & w12049) | (~w12341 & w13639) | (w12049 & w13639);
assign w12343 = ~w12059 & ~w12064;
assign w12344 = w12343 & w14071;
assign w12345 = ~w12058 & w12344;
assign w12346 = ~w12054 & ~w12345;
assign w12347 = ~w12060 & ~w12065;
assign w12348 = (~w12347 & w12054) | (~w12347 & w13640) | (w12054 & w13640);
assign w12349 = ~w12082 & ~w12087;
assign w12350 = w12349 & w14072;
assign w12351 = ~w12081 & w12350;
assign w12352 = ~w12083 & ~w12088;
assign w12353 = (~w12352 & w12077) | (~w12352 & w13641) | (w12077 & w13641);
assign w12354 = ~w12348 & w12353;
assign w12355 = w12348 & ~w12353;
assign w12356 = ~w12354 & ~w12355;
assign w12357 = ~w12342 & ~w12356;
assign w12358 = ~w12341 & w12356;
assign w12359 = ~w12339 & w12358;
assign w12360 = ~w12357 & ~w12359;
assign w12361 = ~w12017 & ~w12040;
assign w12362 = ~w11994 & ~w12361;
assign w12363 = ~w12016 & ~w12039;
assign w12364 = w12363 & w13172;
assign w12365 = (~w12364 & w11994) | (~w12364 & w13642) | (w11994 & w13642);
assign w12366 = ~w12004 & ~w12009;
assign w12367 = w12366 & w14073;
assign w12368 = ~w12003 & w12367;
assign w12369 = ~w11999 & ~w12368;
assign w12370 = ~w12005 & ~w12010;
assign w12371 = (~w12370 & w11999) | (~w12370 & w13643) | (w11999 & w13643);
assign w12372 = ~w12027 & ~w12032;
assign w12373 = w12372 & w14074;
assign w12374 = ~w12026 & w12373;
assign w12375 = ~w12028 & ~w12033;
assign w12376 = (~w12375 & w12022) | (~w12375 & w13644) | (w12022 & w13644);
assign w12377 = ~w12371 & w12376;
assign w12378 = w12371 & ~w12376;
assign w12379 = ~w12377 & ~w12378;
assign w12380 = ~w12365 & ~w12379;
assign w12381 = ~w12364 & w12379;
assign w12382 = ~w12362 & w12381;
assign w12383 = ~w12380 & ~w12382;
assign w12384 = ~w12360 & w12383;
assign w12385 = w12360 & ~w12383;
assign w12386 = ~w12384 & ~w12385;
assign w12387 = ~w12337 & ~w12386;
assign w12388 = w12337 & w12386;
assign w12389 = ~w12387 & ~w12388;
assign w12390 = ~w12334 & w12389;
assign w12391 = w12334 & ~w12389;
assign w12392 = ~w12390 & ~w12391;
assign w12393 = ~w12306 & ~w12392;
assign w12394 = w12306 & w12392;
assign w12395 = ~w12393 & ~w12394;
assign w12396 = ~w12240 & ~w12293;
assign w12397 = w12240 & w12293;
assign w12398 = (~w12397 & w12187) | (~w12397 & w13994) | (w12187 & w13994);
assign w12399 = ~w12265 & ~w12287;
assign w12400 = ~w12243 & ~w12399;
assign w12401 = ~w12264 & ~w12286;
assign w12402 = w12401 & w13995;
assign w12403 = ~w12252 & ~w12257;
assign w12404 = (w12403 & w11827) | (w12403 & w13996) | (w11827 & w13996);
assign w12405 = ~w12251 & w12404;
assign w12406 = (~w12405 & w12245) | (~w12405 & w13997) | (w12245 & w13997);
assign w12407 = ~w12253 & ~w12258;
assign w12408 = (~w12245 & w13998) | (~w12245 & w13999) | (w13998 & w13999);
assign w12409 = ~w12274 & ~w12279;
assign w12410 = (w12409 & w11780) | (w12409 & w14000) | (w11780 & w14000);
assign w12411 = ~w12273 & w12410;
assign w12412 = ~w12275 & ~w12280;
assign w12413 = (~w12267 & w14002) | (~w12267 & w14003) | (w14002 & w14003);
assign w12414 = ~w12408 & w12413;
assign w12415 = w12408 & ~w12413;
assign w12416 = ~w12414 & ~w12415;
assign w12417 = (~w12416 & w12400) | (~w12416 & w14004) | (w12400 & w14004);
assign w12418 = ~w12402 & w12416;
assign w12419 = ~w12400 & w12418;
assign w12420 = ~w12417 & ~w12419;
assign w12421 = ~w12212 & ~w12234;
assign w12422 = ~w12190 & ~w12421;
assign w12423 = ~w12211 & ~w12233;
assign w12424 = w12423 & w14005;
assign w12425 = ~w12199 & ~w12204;
assign w12426 = (w12425 & w11930) | (w12425 & w14006) | (w11930 & w14006);
assign w12427 = ~w12198 & w12426;
assign w12428 = (~w12427 & w12192) | (~w12427 & w14007) | (w12192 & w14007);
assign w12429 = ~w12200 & ~w12205;
assign w12430 = (~w12192 & w14008) | (~w12192 & w14009) | (w14008 & w14009);
assign w12431 = ~w12221 & ~w12226;
assign w12432 = (w12431 & w11883) | (w12431 & w14010) | (w11883 & w14010);
assign w12433 = ~w12220 & w12432;
assign w12434 = ~w12222 & ~w12227;
assign w12435 = (~w12214 & w14012) | (~w12214 & w14013) | (w14012 & w14013);
assign w12436 = ~w12430 & w12435;
assign w12437 = w12430 & ~w12435;
assign w12438 = ~w12436 & ~w12437;
assign w12439 = (~w12438 & w12422) | (~w12438 & w14014) | (w12422 & w14014);
assign w12440 = ~w12424 & w12438;
assign w12441 = ~w12422 & w12440;
assign w12442 = ~w12439 & ~w12441;
assign w12443 = ~w12420 & w12442;
assign w12444 = w12420 & ~w12442;
assign w12445 = ~w12443 & ~w12444;
assign w12446 = ~w12398 & ~w12445;
assign w12447 = w12398 & w12445;
assign w12448 = ~w12446 & ~w12447;
assign w12449 = ~w12395 & ~w12448;
assign w12450 = ~w12393 & w12448;
assign w12451 = ~w12394 & w12450;
assign w12452 = (~w12451 & w12303) | (~w12451 & w13789) | (w12303 & w13789);
assign w12453 = ~w12334 & ~w12389;
assign w12454 = w12334 & w12389;
assign w12455 = (~w12454 & w12306) | (~w12454 & w13790) | (w12306 & w13790);
assign w12456 = ~w12319 & ~w12324;
assign w12457 = (~w12310 & w14015) | (~w12310 & w14016) | (w14015 & w14016);
assign w12458 = ~w12328 & ~w12456;
assign w12459 = (w12458 & w12310) | (w12458 & w13792) | (w12310 & w13792);
assign w12460 = ~w12457 & ~w12459;
assign w12461 = ~w12360 & ~w12383;
assign w12462 = ~w12337 & ~w12461;
assign w12463 = ~w12359 & ~w12382;
assign w12464 = w12463 & w13645;
assign w12465 = (~w12464 & w12337) | (~w12464 & w13793) | (w12337 & w13793);
assign w12466 = ~w12370 & ~w12375;
assign w12467 = (w12466 & w12022) | (w12466 & w14017) | (w12022 & w14017);
assign w12468 = ~w12369 & w12467;
assign w12469 = ~w12365 & ~w12468;
assign w12470 = ~w12371 & ~w12376;
assign w12471 = (~w12470 & w12365) | (~w12470 & w13794) | (w12365 & w13794);
assign w12472 = ~w12347 & ~w12352;
assign w12473 = (w12472 & w12077) | (w12472 & w14018) | (w12077 & w14018);
assign w12474 = ~w12346 & w12473;
assign w12475 = ~w12348 & ~w12353;
assign w12476 = (~w12475 & w12342) | (~w12475 & w13795) | (w12342 & w13795);
assign w12477 = ~w12471 & w12476;
assign w12478 = w12471 & ~w12476;
assign w12479 = ~w12477 & ~w12478;
assign w12480 = ~w12465 & ~w12479;
assign w12481 = ~w12464 & w12479;
assign w12482 = ~w12462 & w12481;
assign w12483 = ~w12480 & ~w12482;
assign w12484 = ~w12460 & ~w12483;
assign w12485 = ~w12459 & ~w12482;
assign w12486 = w12485 & w13796;
assign w12487 = ~w12484 & ~w12486;
assign w12488 = ~w12455 & w12487;
assign w12489 = w12455 & ~w12487;
assign w12490 = ~w12488 & ~w12489;
assign w12491 = ~w12420 & ~w12442;
assign w12492 = ~w12398 & ~w12491;
assign w12493 = ~w12419 & ~w12441;
assign w12494 = w12493 & w14019;
assign w12495 = ~w12429 & ~w12434;
assign w12496 = w12495 & w14075;
assign w12497 = ~w12428 & w12496;
assign w12498 = (~w12497 & w12422) | (~w12497 & w14020) | (w12422 & w14020);
assign w12499 = ~w12430 & ~w12435;
assign w12500 = (~w12422 & w14021) | (~w12422 & w14022) | (w14021 & w14022);
assign w12501 = ~w12407 & ~w12412;
assign w12502 = w12501 & w14076;
assign w12503 = ~w12406 & w12502;
assign w12504 = ~w12408 & ~w12413;
assign w12505 = (~w12400 & w14024) | (~w12400 & w14025) | (w14024 & w14025);
assign w12506 = ~w12500 & w12505;
assign w12507 = w12500 & ~w12505;
assign w12508 = ~w12506 & ~w12507;
assign w12509 = (~w12508 & w12492) | (~w12508 & w14026) | (w12492 & w14026);
assign w12510 = ~w12494 & w12508;
assign w12511 = ~w12492 & w12510;
assign w12512 = ~w12509 & ~w12511;
assign w12513 = ~w12490 & ~w12512;
assign w12514 = ~w12452 & ~w12513;
assign w12515 = ~w12488 & w12512;
assign w12516 = ~w12489 & w12515;
assign w12517 = (~w12516 & w12452) | (~w12516 & w14027) | (w12452 & w14027);
assign w12518 = ~w12455 & ~w12484;
assign w12519 = (~w12486 & w12455) | (~w12486 & w14028) | (w12455 & w14028);
assign w12520 = ~w12470 & ~w12475;
assign w12521 = (w12520 & w12342) | (w12520 & w14029) | (w12342 & w14029);
assign w12522 = ~w12469 & w12521;
assign w12523 = ~w12465 & ~w12522;
assign w12524 = ~w12471 & ~w12476;
assign w12525 = ~w12457 & ~w12524;
assign w12526 = ~w12523 & w12525;
assign w12527 = (~w12524 & w12465) | (~w12524 & w14030) | (w12465 & w14030);
assign w12528 = w12457 & ~w12527;
assign w12529 = ~w12526 & ~w12528;
assign w12530 = ~w12519 & w12529;
assign w12531 = ~w12486 & ~w12529;
assign w12532 = ~w12518 & w12531;
assign w12533 = ~w12530 & ~w12532;
assign w12534 = ~w12499 & ~w12504;
assign w12535 = w12534 & w14077;
assign w12536 = ~w12498 & w12535;
assign w12537 = ~w12500 & ~w12505;
assign w12538 = (~w12492 & w14031) | (~w12492 & w14032) | (w14031 & w14032);
assign w12539 = ~w12533 & w12538;
assign w12540 = (~w12538 & w12518) | (~w12538 & w14033) | (w12518 & w14033);
assign w12541 = ~w12530 & w12540;
assign w12542 = (~w12541 & w12517) | (~w12541 & w14034) | (w12517 & w14034);
assign w12543 = (~w12528 & w12519) | (~w12528 & w14035) | (w12519 & w14035);
assign w12544 = ~w12542 & w12543;
assign w12545 = ~w12541 & ~w12543;
assign w12546 = (w12545 & w12517) | (w12545 & w14036) | (w12517 & w14036);
assign w12547 = ~w12544 & ~w12546;
assign w12548 = ~w12533 & ~w12538;
assign w12549 = (w12538 & w12518) | (w12538 & w14037) | (w12518 & w14037);
assign w12550 = ~w12530 & w12549;
assign w12551 = ~w12516 & ~w12550;
assign w12552 = ~w12514 & w14038;
assign w12553 = ~w12548 & ~w12550;
assign w12554 = ~w12517 & ~w12553;
assign w12555 = ~w12490 & w12512;
assign w12556 = ~w12488 & ~w12512;
assign w12557 = ~w12489 & w12556;
assign w12558 = ~w12555 & ~w12557;
assign w12559 = w12452 & w12558;
assign w12560 = ~w12452 & ~w12558;
assign w12561 = ~w12393 & ~w12448;
assign w12562 = ~w12394 & w12561;
assign w12563 = ~w12395 & w12448;
assign w12564 = ~w12562 & ~w12563;
assign w12565 = w12303 & w12564;
assign w12566 = ~w12303 & ~w12564;
assign w12567 = ~w12184 & w12299;
assign w12568 = ~w12182 & ~w12299;
assign w12569 = ~w12183 & w12568;
assign w12570 = ~w12567 & ~w12569;
assign w12571 = w11985 & w12570;
assign w12572 = ~w11985 & ~w12570;
assign w12573 = ~w11764 & ~w11981;
assign w12574 = ~w11765 & w12573;
assign w12575 = ~w11766 & w11981;
assign w12576 = ~w12574 & ~w12575;
assign w12577 = w11416 & w12576;
assign w12578 = ~w11416 & ~w12576;
assign w12579 = ~w10894 & w11412;
assign w12580 = (~w11412 & w10891) | (~w11412 & w14039) | (w10891 & w14039);
assign w12581 = ~w10893 & w12580;
assign w12582 = ~w12579 & ~w12581;
assign w12583 = w10075 & w12582;
assign w12584 = ~w10075 & ~w12582;
assign w12585 = (~w10071 & w9372) | (~w10071 & w12953) | (w9372 & w12953);
assign w12586 = ~w9374 & w12585;
assign w12587 = ~w9375 & w10071;
assign w12588 = (~w8254 & w12587) | (~w8254 & w14040) | (w12587 & w14040);
assign w12589 = ~w8240 & ~w8241;
assign w12590 = ~w8242 & w12589;
assign w12591 = w8240 & ~w8243;
assign w12592 = ~w12590 & ~w12591;
assign w12593 = A_1000 & ~w12592;
assign w12594 = (~w12587 & w14041) | (~w12587 & w14042) | (w14041 & w14042);
assign w12595 = ~w12587 & w13474;
assign w12596 = w8244 & ~w8248;
assign w12597 = ~w8237 & w12596;
assign w12598 = ~w8244 & ~w8252;
assign w12599 = ~w12597 & ~w12598;
assign w12600 = w3162 & ~w12599;
assign w12601 = ~w8250 & ~w8253;
assign w12602 = ~w3162 & ~w12601;
assign w12603 = ~w12600 & ~w12602;
assign w12604 = ~w12595 & ~w12603;
assign w12605 = w12594 & w12604;
assign w12606 = w12605 & w12621;
assign w12607 = w12606 & w12632;
assign w12608 = w12607 & w12636;
assign w12609 = w12608 & w12619;
assign w12610 = w12609 & w12617;
assign w12611 = w12610 & w12615;
assign w12612 = w12547 & w12611;
assign w12613 = ~w12547 & ~w12611;
assign w12614 = ~w12612 & ~w12613;
assign w12615 = ~w12552 & ~w12554;
assign w12616 = ~w12610 & ~w12615;
assign w12617 = ~w12559 & ~w12560;
assign w12618 = ~w12609 & ~w12617;
assign w12619 = ~w12565 & ~w12566;
assign w12620 = ~w12608 & ~w12619;
assign w12621 = ~w12583 & ~w12584;
assign w12622 = ~w12605 & ~w12621;
assign w12623 = w12593 & ~w12603;
assign w12624 = (~w12623 & w12588) | (~w12623 & w13475) | (w12588 & w13475);
assign w12625 = ~w12605 & ~w12624;
assign w12626 = (w12593 & w12599) | (w12593 & w14043) | (w12599 & w14043);
assign w12627 = ~w12602 & w12626;
assign w12628 = ~w12593 & ~w12603;
assign w12629 = ~w12627 & ~w12628;
assign w12630 = ~w12625 & w12629;
assign w12631 = ~w12630 & w12657;
assign w12632 = ~w12577 & ~w12578;
assign w12633 = ~w12606 & ~w12632;
assign w12634 = ~w12607 & ~w12633;
assign w12635 = ~w12631 & ~w12634;
assign w12636 = ~w12571 & ~w12572;
assign w12637 = ~w12607 & ~w12636;
assign w12638 = ~w12608 & ~w12637;
assign w12639 = ~w12635 & w12638;
assign w12640 = w12639 & w12681;
assign w12641 = w12640 & w12656;
assign w12642 = w12641 & w12690;
assign w12643 = ~w12614 & w12642;
assign w12644 = ~w12547 & w12611;
assign w12645 = ~w12542 & ~w12543;
assign w12646 = ~w12644 & w12645;
assign w12647 = w12611 & ~w12645;
assign w12648 = ~w12547 & w12647;
assign w12649 = ~w12543 & w12609;
assign w12650 = w12617 & w12649;
assign w12651 = w12650 & w14044;
assign w12652 = ~w12547 & w12651;
assign w12653 = ~w12648 & ~w12652;
assign w12654 = ~w12646 & w12653;
assign w12655 = ~w12643 & w12654;
assign w12656 = ~w12610 & ~w12618;
assign w12657 = ~w12606 & ~w12622;
assign w12658 = w12630 & ~w12657;
assign w12659 = ~w12631 & ~w12658;
assign w12660 = w12625 & ~w12629;
assign w12661 = (A_1000 & ~w12589) | (A_1000 & w14045) | (~w12589 & w14045);
assign w12662 = ~w12591 & w12661;
assign w12663 = ~A_1000 & ~w12592;
assign w12664 = ~w12662 & ~w12663;
assign w12665 = (w12664 & w12625) | (w12664 & w12954) | (w12625 & w12954);
assign w12666 = ~w12660 & w12665;
assign w12667 = w12625 & ~w12666;
assign w12668 = ~w12630 & ~w12660;
assign w12669 = ~w12664 & ~w12668;
assign w12670 = ~w12667 & ~w12669;
assign w12671 = (w12657 & ~w12670) | (w12657 & w13173) | (~w12670 & w13173);
assign w12672 = (~w12631 & w12671) | (~w12631 & w12955) | (w12671 & w12955);
assign w12673 = w12631 & w12634;
assign w12674 = w12635 & ~w12638;
assign w12675 = ~w12639 & ~w12674;
assign w12676 = ~w12673 & ~w12675;
assign w12677 = (w12638 & ~w12676) | (w12638 & w12956) | (~w12676 & w12956);
assign w12678 = (~w12955 & w13174) | (~w12955 & w13175) | (w13174 & w13175);
assign w12679 = (~w13175 & w13476) | (~w13175 & w13477) | (w13476 & w13477);
assign w12680 = (w12639 & w12677) | (w12639 & w13176) | (w12677 & w13176);
assign w12681 = ~w12609 & ~w12620;
assign w12682 = ~w12639 & w12681;
assign w12683 = ~w12640 & ~w12656;
assign w12684 = ~w12641 & ~w12683;
assign w12685 = ~w12682 & ~w12684;
assign w12686 = (w12656 & ~w12685) | (w12656 & w12957) | (~w12685 & w12957);
assign w12687 = w12641 & ~w12642;
assign w12688 = (w12687 & w12686) | (w12687 & w13647) | (w12686 & w13647);
assign w12689 = w12642 & ~w12686;
assign w12690 = ~w12611 & ~w12616;
assign w12691 = (w12690 & ~w12689) | (w12690 & w12958) | (~w12689 & w12958);
assign w12692 = w12642 & ~w12643;
assign w12693 = (w12692 & w12691) | (w12692 & w13648) | (w12691 & w13648);
assign w12694 = w12643 & ~w12688;
assign w12695 = (w12694 & w13177) | (w12694 & w13178) | (w13177 & w13178);
assign w12696 = w12642 & ~w12648;
assign w12697 = w12696 & w14046;
assign w12698 = ~w12646 & ~w12648;
assign w12699 = ~w12643 & w12698;
assign w12700 = w12652 & ~w12699;
assign w12701 = (~w12697 & w12700) | (~w12697 & w13179) | (w12700 & w13179);
assign w12702 = (w12701 & ~w12695) | (w12701 & w13649) | (~w12695 & w13649);
assign w12703 = w12655 & ~w12702;
assign w12704 = ~A_18 & ~w3577;
assign w12705 = ~A_15 & ~w3582;
assign w12706 = ~A_30 & ~w3659;
assign w12707 = ~A_27 & ~w3664;
assign w12708 = ~A_48 & ~w3843;
assign w12709 = ~A_45 & ~w3848;
assign w12710 = ~A_54 & ~w3877;
assign w12711 = ~A_51 & ~w3882;
assign w12712 = ~A_42 & ~w3946;
assign w12713 = ~A_39 & ~w3948;
assign w12714 = ~A_36 & ~w3979;
assign w12715 = ~A_33 & ~w3981;
assign w12716 = ~A_60 & ~w4026;
assign w12717 = ~A_57 & ~w4031;
assign w12718 = ~A_66 & ~w4060;
assign w12719 = ~A_63 & ~w4065;
assign w12720 = ~A_72 & ~w4108;
assign w12721 = ~A_69 & ~w4113;
assign w12722 = ~A_78 & ~w4142;
assign w12723 = ~A_75 & ~w4147;
assign w12724 = ~A_204 & ~w5057;
assign w12725 = ~A_201 & ~w5062;
assign w12726 = ~A_210 & ~w5091;
assign w12727 = ~A_207 & ~w5096;
assign w12728 = ~A_216 & ~w5139;
assign w12729 = ~A_213 & ~w5144;
assign w12730 = ~A_222 & ~w5173;
assign w12731 = ~A_219 & ~w5178;
assign w12732 = ~A_198 & ~w5258;
assign w12733 = ~A_195 & ~w5260;
assign w12734 = ~A_192 & ~w5291;
assign w12735 = ~A_189 & ~w5293;
assign w12736 = ~A_186 & ~w5327;
assign w12737 = ~A_183 & ~w5329;
assign w12738 = ~A_180 & ~w5360;
assign w12739 = ~A_177 & ~w5362;
assign w12740 = ~A_240 & ~w5438;
assign w12741 = ~A_237 & ~w5443;
assign w12742 = ~A_246 & ~w5472;
assign w12743 = ~A_243 & ~w5477;
assign w12744 = ~A_234 & ~w5541;
assign w12745 = ~A_231 & ~w5543;
assign w12746 = ~A_228 & ~w5574;
assign w12747 = ~A_225 & ~w5576;
assign w12748 = ~A_252 & ~w5621;
assign w12749 = ~A_249 & ~w5626;
assign w12750 = ~A_258 & ~w5655;
assign w12751 = ~A_255 & ~w5660;
assign w12752 = ~A_264 & ~w5703;
assign w12753 = ~A_261 & ~w5708;
assign w12754 = ~A_270 & ~w5737;
assign w12755 = ~A_267 & ~w5742;
assign w12756 = ~A_174 & ~w5856;
assign w12757 = ~A_171 & ~w5858;
assign w12758 = ~A_168 & ~w5889;
assign w12759 = ~A_165 & ~w5891;
assign w12760 = ~A_162 & ~w5925;
assign w12761 = ~A_159 & ~w5927;
assign w12762 = ~A_156 & ~w5958;
assign w12763 = ~A_153 & ~w5960;
assign w12764 = ~A_150 & ~w5997;
assign w12765 = ~A_147 & ~w5999;
assign w12766 = ~A_144 & ~w6030;
assign w12767 = ~A_141 & ~w6032;
assign w12768 = ~A_138 & ~w6066;
assign w12769 = ~A_135 & ~w6068;
assign w12770 = ~A_132 & ~w6099;
assign w12771 = ~A_129 & ~w6101;
assign w12772 = ~A_126 & ~w6141;
assign w12773 = ~A_123 & ~w6143;
assign w12774 = ~A_120 & ~w6174;
assign w12775 = ~A_117 & ~w6176;
assign w12776 = ~A_114 & ~w6210;
assign w12777 = ~A_111 & ~w6212;
assign w12778 = ~A_108 & ~w6243;
assign w12779 = ~A_105 & ~w6245;
assign w12780 = ~A_102 & ~w6282;
assign w12781 = ~A_99 & ~w6284;
assign w12782 = ~A_96 & ~w6315;
assign w12783 = ~A_93 & ~w6317;
assign w12784 = ~A_90 & ~w6351;
assign w12785 = ~A_87 & ~w6353;
assign w12786 = ~A_84 & ~w6384;
assign w12787 = ~A_81 & ~w6386;
assign w12788 = ~A_336 & ~w6633;
assign w12789 = ~A_333 & ~w6638;
assign w12790 = ~A_342 & ~w6667;
assign w12791 = ~A_339 & ~w6672;
assign w12792 = ~A_330 & ~w6736;
assign w12793 = ~A_327 & ~w6738;
assign w12794 = ~A_324 & ~w6769;
assign w12795 = ~A_321 & ~w6771;
assign w12796 = ~A_348 & ~w6816;
assign w12797 = ~A_345 & ~w6821;
assign w12798 = ~A_354 & ~w6850;
assign w12799 = ~A_351 & ~w6855;
assign w12800 = ~A_360 & ~w6898;
assign w12801 = ~A_357 & ~w6903;
assign w12802 = ~A_366 & ~w6932;
assign w12803 = ~A_363 & ~w6937;
assign w12804 = ~A_318 & ~w7034;
assign w12805 = ~A_315 & ~w7036;
assign w12806 = ~A_312 & ~w7067;
assign w12807 = ~A_309 & ~w7069;
assign w12808 = ~A_306 & ~w7103;
assign w12809 = ~A_303 & ~w7105;
assign w12810 = ~A_300 & ~w7136;
assign w12811 = ~A_297 & ~w7138;
assign w12812 = ~A_294 & ~w7175;
assign w12813 = ~A_291 & ~w7177;
assign w12814 = ~A_288 & ~w7208;
assign w12815 = ~A_285 & ~w7210;
assign w12816 = ~A_282 & ~w7244;
assign w12817 = ~A_279 & ~w7246;
assign w12818 = ~A_276 & ~w7277;
assign w12819 = ~A_273 & ~w7279;
assign w12820 = ~A_396 & ~w7413;
assign w12821 = ~A_393 & ~w7418;
assign w12822 = ~A_402 & ~w7447;
assign w12823 = ~A_399 & ~w7452;
assign w12824 = ~A_408 & ~w7495;
assign w12825 = ~A_405 & ~w7500;
assign w12826 = ~A_414 & ~w7529;
assign w12827 = ~A_411 & ~w7534;
assign w12828 = ~A_390 & ~w7614;
assign w12829 = ~A_387 & ~w7616;
assign w12830 = ~A_384 & ~w7647;
assign w12831 = ~A_381 & ~w7649;
assign w12832 = ~A_378 & ~w7683;
assign w12833 = ~A_375 & ~w7685;
assign w12834 = ~A_372 & ~w7716;
assign w12835 = ~A_369 & ~w7718;
assign w12836 = ~A_432 & ~w7794;
assign w12837 = ~A_429 & ~w7799;
assign w12838 = ~A_438 & ~w7828;
assign w12839 = ~A_435 & ~w7833;
assign w12840 = ~A_426 & ~w7897;
assign w12841 = ~A_423 & ~w7899;
assign w12842 = ~A_420 & ~w7930;
assign w12843 = ~A_417 & ~w7932;
assign w12844 = ~A_444 & ~w7976;
assign w12845 = ~A_441 & ~w7981;
assign w12846 = ~A_450 & ~w8010;
assign w12847 = ~A_447 & ~w8015;
assign w12848 = ~A_456 & ~w8058;
assign w12849 = ~A_453 & ~w8063;
assign w12850 = ~A_462 & ~w8092;
assign w12851 = ~A_459 & ~w8097;
assign w12852 = w8133 & w8090;
assign w12853 = ~w8149 & ~w8134;
assign w12854 = w8134 & w8149;
assign w12855 = w8149 & ~w8134;
assign w12856 = w8154 & w8057;
assign w12857 = ~w4253 & w12959;
assign w12858 = ~w4235 & w12960;
assign w12859 = w3820 & w12961;
assign w12860 = (w12962 & w3777) | (w12962 & w13180) | (w3777 & w13180);
assign w12861 = w8267 & w8275;
assign w12862 = ~w8265 & ~w8279;
assign w12863 = w4008 & w4003;
assign w12864 = w3913 & w3875;
assign w12865 = w4096 & w4058;
assign w12866 = w4178 & w4140;
assign w12867 = w8260 & ~w8666;
assign w12868 = w6596 & w6591;
assign w12869 = w6575 & w6570;
assign w12870 = w6527 & w6522;
assign w12871 = w6545 & w6540;
assign w12872 = w6444 & w6439;
assign w12873 = w6423 & w6418;
assign w12874 = w6468 & w6463;
assign w12875 = w6486 & w6481;
assign w12876 = w5414 & w5409;
assign w12877 = w5393 & w5388;
assign w12878 = w5127 & w5089;
assign w12879 = w5209 & w5171;
assign w12880 = w5603 & w5598;
assign w12881 = w5508 & w5470;
assign w12882 = w5691 & w5653;
assign w12883 = w5773 & w5735;
assign w12884 = w7382 & w7377;
assign w12885 = w7361 & w7356;
assign w12886 = w7313 & w7308;
assign w12887 = w7331 & w7326;
assign w12888 = w6798 & w6793;
assign w12889 = w6703 & w6665;
assign w12890 = w6886 & w6848;
assign w12891 = w6968 & w6930;
assign w12892 = w7770 & w7765;
assign w12893 = w7749 & w7744;
assign w12894 = w7483 & w7445;
assign w12895 = w7565 & w7527;
assign w12896 = w7959 & w7954;
assign w12897 = w7864 & w7826;
assign w12898 = w8046 & w8008;
assign w12899 = w8128 & w8090;
assign w12900 = ~w9335 & ~w9321;
assign w12901 = w7973 & ~w10118;
assign w12902 = ~w9299 & ~w9285;
assign w12903 = w10147 & ~w10148;
assign w12904 = w7588 & ~w10150;
assign w12905 = ~w9255 & ~w9241;
assign w12906 = w7784 & ~w10173;
assign w12907 = ~w9219 & ~w9205;
assign w12908 = w10208 & ~w10209;
assign w12909 = w10211 & ~w10212;
assign w12910 = w6991 & ~w10214;
assign w12911 = ~w9167 & ~w9153;
assign w12912 = w6812 & ~w10237;
assign w12913 = ~w9131 & ~w9117;
assign w12914 = w10266 & ~w10267;
assign w12915 = w7344 & ~w10269;
assign w12916 = ~w9087 & ~w9073;
assign w12917 = w7396 & ~w10292;
assign w12918 = ~w9051 & ~w9037;
assign w12919 = w10333 & ~w10334;
assign w12920 = w10336 & ~w10337;
assign w12921 = w10339 & ~w10340;
assign w12922 = w5796 & ~w10342;
assign w12923 = ~w8991 & ~w8977;
assign w12924 = w5617 & ~w10365;
assign w12925 = ~w8955 & ~w8941;
assign w12926 = w10394 & ~w10395;
assign w12927 = w5232 & ~w10397;
assign w12928 = ~w8911 & ~w8897;
assign w12929 = w5428 & ~w10420;
assign w12930 = ~w8875 & ~w8861;
assign w12931 = w10455 & ~w10456;
assign w12932 = w10458 & ~w10459;
assign w12933 = w6499 & ~w10461;
assign w12934 = ~w8823 & ~w8809;
assign w12935 = w6458 & ~w10484;
assign w12936 = ~w8787 & ~w8773;
assign w12937 = w10513 & ~w10514;
assign w12938 = w6558 & ~w10516;
assign w12939 = ~w8743 & ~w8729;
assign w12940 = w6610 & ~w10539;
assign w12941 = ~w8707 & ~w8693;
assign w12942 = w10595 & ~w10596;
assign w12943 = w10598 & ~w10599;
assign w12944 = w4201 & ~w10601;
assign w12945 = ~w8390 & ~w8376;
assign w12946 = w4022 & ~w10624;
assign w12947 = ~w8354 & ~w8340;
assign w12948 = w10653 & ~w10655;
assign w12949 = w8275 & w8265;
assign w12950 = ~w8310 & ~w8296;
assign w12951 = w10669 & ~w10682;
assign w12952 = w10669 & ~w11433;
assign w12953 = w8256 & ~w10071;
assign w12954 = (w12664 & w12628) | (w12664 & w14047) | (w12628 & w14047);
assign w12955 = ~w12670 & w13181;
assign w12956 = w12672 & w12638;
assign w12957 = (w12963 & w12677) | (w12963 & w13650) | (w12677 & w13650);
assign w12958 = (w12964 & w12680) | (w12964 & w14048) | (w12680 & w14048);
assign w12959 = ~w3542 & ~w5049;
assign w12960 = ~w3842 & ~w3542;
assign w12961 = ~w3816 & w3801;
assign w12962 = ~w3786 & ~w3818;
assign w12963 = w12639 & w12656;
assign w12964 = w12684 & w12690;
assign w12965 = ~w12614 & w12690;
assign w12966 = (w12680 & w14066) | (w12680 & w14067) | (w14066 & w14067);
assign w12967 = ~A_12 & ~w3543;
assign w12968 = ~A_9 & ~w3548;
assign w12969 = ~A_24 & ~w3625;
assign w12970 = ~A_21 & ~w3630;
assign w12971 = w3700 & w3657;
assign w12972 = ~w3716 & ~w3701;
assign w12973 = w3716 & ~w3701;
assign w12974 = w3721 & w3624;
assign w12975 = w3768 & A_6;
assign w12976 = w3774 & ~w3766;
assign w12977 = w3918 & w3875;
assign w12978 = ~w3998 & ~w3919;
assign w12979 = w4183 & w4140;
assign w12980 = ~w4199 & ~w4184;
assign w12981 = w4184 & w4199;
assign w12982 = w4199 & ~w4184;
assign w12983 = w4204 & w4107;
assign w12984 = w5214 & w5171;
assign w12985 = ~w5230 & ~w5215;
assign w12986 = w5215 & w5230;
assign w12987 = w5230 & ~w5215;
assign w12988 = w5235 & w5138;
assign w12989 = w5398 & w5388;
assign w12990 = ~w5404 & ~w5399;
assign w12991 = w5513 & w5470;
assign w12992 = ~w5593 & ~w5514;
assign w12993 = w5778 & w5735;
assign w12994 = ~w5794 & ~w5779;
assign w12995 = w5779 & w5794;
assign w12996 = w5794 & ~w5779;
assign w12997 = w5799 & w5702;
assign w12998 = w6428 & w6418;
assign w12999 = ~w6434 & ~w6429;
assign w13000 = w6491 & w6481;
assign w13001 = ~w6497 & ~w6492;
assign w13002 = w6492 & w6497;
assign w13003 = w6497 & ~w6492;
assign w13004 = w6502 & w6479;
assign w13005 = w6550 & w6540;
assign w13006 = ~w6556 & ~w6551;
assign w13007 = w6551 & w6556;
assign w13008 = w6556 & ~w6551;
assign w13009 = w6561 & w6538;
assign w13010 = w6580 & w6570;
assign w13011 = ~w6586 & ~w6581;
assign w13012 = w6708 & w6665;
assign w13013 = ~w6788 & ~w6709;
assign w13014 = w6973 & w6930;
assign w13015 = ~w6989 & ~w6974;
assign w13016 = w6974 & w6989;
assign w13017 = w6989 & ~w6974;
assign w13018 = w6994 & w6897;
assign w13019 = w7336 & w7326;
assign w13020 = ~w7342 & ~w7337;
assign w13021 = w7337 & w7342;
assign w13022 = w7342 & ~w7337;
assign w13023 = w7347 & w7324;
assign w13024 = w7366 & w7356;
assign w13025 = ~w7372 & ~w7367;
assign w13026 = w7570 & w7527;
assign w13027 = ~w7586 & ~w7571;
assign w13028 = w7571 & w7586;
assign w13029 = w7586 & ~w7571;
assign w13030 = w7591 & w7494;
assign w13031 = w7754 & w7744;
assign w13032 = ~w7760 & ~w7755;
assign w13033 = w7869 & w7826;
assign w13034 = w7949 & ~w7870;
assign w13035 = w7870 & ~w7949;
assign w13036 = ~w7949 & ~w7870;
assign w13037 = w7972 & ~w7970;
assign w13038 = w8055 & w8008;
assign w13039 = w8134 & ~w8149;
assign w13040 = ~w8163 & ~w8057;
assign w13041 = ~w8163 & ~w8155;
assign w13042 = w8165 & ~w7975;
assign w13043 = ~w7975 & ~w8180;
assign w13044 = w8168 & w8180;
assign w13045 = ~w7975 & w8180;
assign w13046 = w8168 & ~w8180;
assign w13047 = w3613 & w3575;
assign w13048 = w3695 & w3657;
assign w13049 = w10095 & ~w10098;
assign w13050 = w8133 & w9329;
assign w13051 = w8055 & w9315;
assign w13052 = ~w10121 & w10118;
assign w13053 = ~w10121 & ~w9274;
assign w13054 = w7869 & w9293;
assign w13055 = w7968 & w9279;
assign w13056 = ~w10153 & w10150;
assign w13057 = ~w10153 & ~w9230;
assign w13058 = w7570 & w9249;
assign w13059 = w7492 & w9235;
assign w13060 = ~w10176 & w10173;
assign w13061 = ~w10176 & ~w9194;
assign w13062 = w7754 & w9213;
assign w13063 = w7779 & w9199;
assign w13064 = ~w10217 & w10214;
assign w13065 = ~w10217 & ~w9142;
assign w13066 = w6973 & w9161;
assign w13067 = w6895 & w9147;
assign w13068 = ~w10240 & w10237;
assign w13069 = ~w10240 & ~w9106;
assign w13070 = w6708 & w9125;
assign w13071 = w6807 & w9111;
assign w13072 = ~w10272 & w10269;
assign w13073 = ~w10272 & ~w9062;
assign w13074 = w7336 & w9081;
assign w13075 = w7322 & w9067;
assign w13076 = ~w10295 & w10292;
assign w13077 = ~w10295 & ~w9026;
assign w13078 = w7366 & w9045;
assign w13079 = w7391 & w9031;
assign w13080 = ~w10345 & w10342;
assign w13081 = ~w10345 & ~w8966;
assign w13082 = w5778 & w8985;
assign w13083 = w5700 & w8971;
assign w13084 = ~w10368 & w10365;
assign w13085 = ~w10368 & ~w8930;
assign w13086 = w5513 & w8949;
assign w13087 = w5612 & w8935;
assign w13088 = ~w10400 & w10397;
assign w13089 = ~w10400 & ~w8886;
assign w13090 = w5214 & w8905;
assign w13091 = w5136 & w8891;
assign w13092 = ~w10423 & w10420;
assign w13093 = ~w10423 & ~w8850;
assign w13094 = w5398 & w8869;
assign w13095 = w5423 & w8855;
assign w13096 = ~w10464 & w10461;
assign w13097 = ~w10464 & ~w8798;
assign w13098 = w6491 & w8817;
assign w13099 = w6477 & w8803;
assign w13100 = ~w10487 & w10484;
assign w13101 = ~w10487 & ~w8762;
assign w13102 = w6428 & w8781;
assign w13103 = w6453 & w8767;
assign w13104 = ~w10519 & w10516;
assign w13105 = ~w10519 & ~w8718;
assign w13106 = w6550 & w8737;
assign w13107 = w6536 & w8723;
assign w13108 = ~w10542 & w10539;
assign w13109 = ~w10542 & ~w8682;
assign w13110 = w6580 & w8701;
assign w13111 = w6605 & w8687;
assign w13112 = ~w10604 & w10601;
assign w13113 = ~w10604 & ~w8365;
assign w13114 = w4183 & w8384;
assign w13115 = w4105 & w8370;
assign w13116 = ~w10627 & w10624;
assign w13117 = ~w10627 & ~w8329;
assign w13118 = w3918 & w8348;
assign w13119 = w4017 & w8334;
assign w13120 = ~w10642 & ~w10619;
assign w13121 = ~w10557 & ~w10534;
assign w13122 = ~w10502 & ~w10479;
assign w13123 = ~w10438 & ~w10415;
assign w13124 = ~w10383 & ~w10360;
assign w13125 = ~w10310 & ~w10287;
assign w13126 = ~w10255 & ~w10232;
assign w13127 = ~w10191 & ~w10168;
assign w13128 = ~w10136 & ~w10113;
assign w13129 = w11729 & ~w11731;
assign w13130 = w11733 & ~w11734;
assign w13131 = w11728 & ~w11738;
assign w13132 = w11767 & ~w11768;
assign w13133 = w11770 & ~w11771;
assign w13134 = w11773 & ~w11774;
assign w13135 = w11776 & ~w11779;
assign w13136 = w11795 & ~w11798;
assign w13137 = w11820 & ~w11821;
assign w13138 = w11823 & ~w11826;
assign w13139 = w11842 & ~w11845;
assign w13140 = w11873 & ~w11874;
assign w13141 = w11876 & ~w11877;
assign w13142 = w11879 & ~w11882;
assign w13143 = w11898 & ~w11901;
assign w13144 = w11923 & ~w11924;
assign w13145 = w11926 & ~w11929;
assign w13146 = w11945 & ~w11948;
assign w13147 = w11982 & ~w11984;
assign w13148 = w11986 & ~w11987;
assign w13149 = w11989 & ~w11990;
assign w13150 = w11992 & ~w11993;
assign w13151 = w11995 & ~w11998;
assign w13152 = w11728 & ~w12002;
assign w13153 = w11709 & ~w12008;
assign w13154 = w12018 & ~w12021;
assign w13155 = w11681 & ~w12025;
assign w13156 = w11662 & ~w12031;
assign w13157 = w12047 & ~w12048;
assign w13158 = w12050 & ~w12053;
assign w13159 = w11625 & ~w12057;
assign w13160 = w11606 & ~w12063;
assign w13161 = w12073 & ~w12076;
assign w13162 = w11578 & ~w12080;
assign w13163 = w11559 & ~w12086;
assign w13164 = w12108 & ~w12110;
assign w13165 = w12112 & ~w12115;
assign w13166 = w12117 & ~w12120;
assign w13167 = w11448 & ~w12124;
assign w13168 = w10689 & ~w11437;
assign w13169 = w12149 & ~w12152;
assign w13170 = w12145 & w12171;
assign w13171 = ~w12092 & ~w12069;
assign w13172 = ~w12037 & ~w12014;
assign w13173 = w12659 & w12657;
assign w13174 = ~w12673 & w12631;
assign w13175 = ~w12673 & ~w12671;
assign w13176 = ~w12678 & w13182;
assign w13177 = ~w12643 & w12614;
assign w13178 = (~w12966 & w13651) | (~w12966 & w13652) | (w13651 & w13652);
assign w13179 = w12655 & ~w12697;
assign w13180 = w3779 & w12962;
assign w13181 = w12659 & ~w12631;
assign w13182 = w12675 & w12639;
assign w13183 = ~A_720 & ~w0;
assign w13184 = ~A_717 & ~w5;
assign w13185 = ~A_726 & ~w34;
assign w13186 = ~A_723 & ~w39;
assign w13187 = ~A_714 & ~w103;
assign w13188 = ~A_711 & ~w105;
assign w13189 = ~A_708 & ~w136;
assign w13190 = ~A_705 & ~w138;
assign w13191 = ~A_732 & ~w182;
assign w13192 = ~A_729 & ~w187;
assign w13193 = ~A_738 & ~w216;
assign w13194 = ~A_735 & ~w221;
assign w13195 = ~A_744 & ~w264;
assign w13196 = ~A_741 & ~w269;
assign w13197 = ~A_750 & ~w298;
assign w13198 = ~A_747 & ~w303;
assign w13199 = ~A_702 & ~w399;
assign w13200 = ~A_699 & ~w401;
assign w13201 = ~A_696 & ~w432;
assign w13202 = ~A_693 & ~w434;
assign w13203 = ~A_690 & ~w468;
assign w13204 = ~A_687 & ~w470;
assign w13205 = ~A_684 & ~w501;
assign w13206 = ~A_681 & ~w503;
assign w13207 = ~A_678 & ~w540;
assign w13208 = ~A_675 & ~w542;
assign w13209 = ~A_672 & ~w573;
assign w13210 = ~A_669 & ~w575;
assign w13211 = ~A_666 & ~w609;
assign w13212 = ~A_663 & ~w611;
assign w13213 = ~A_660 & ~w642;
assign w13214 = ~A_657 & ~w644;
assign w13215 = ~A_780 & ~w778;
assign w13216 = ~A_777 & ~w783;
assign w13217 = ~A_786 & ~w812;
assign w13218 = ~A_783 & ~w817;
assign w13219 = ~A_792 & ~w860;
assign w13220 = ~A_789 & ~w865;
assign w13221 = ~A_798 & ~w894;
assign w13222 = ~A_795 & ~w899;
assign w13223 = ~A_774 & ~w979;
assign w13224 = ~A_771 & ~w981;
assign w13225 = ~A_768 & ~w1012;
assign w13226 = ~A_765 & ~w1014;
assign w13227 = ~A_762 & ~w1048;
assign w13228 = ~A_759 & ~w1050;
assign w13229 = ~A_756 & ~w1081;
assign w13230 = ~A_753 & ~w1083;
assign w13231 = ~A_816 & ~w1158;
assign w13232 = ~A_813 & ~w1163;
assign w13233 = ~A_822 & ~w1192;
assign w13234 = ~A_819 & ~w1197;
assign w13235 = ~A_810 & ~w1261;
assign w13236 = ~A_807 & ~w1263;
assign w13237 = ~A_804 & ~w1294;
assign w13238 = ~A_801 & ~w1296;
assign w13239 = ~A_828 & ~w1340;
assign w13240 = ~A_825 & ~w1345;
assign w13241 = ~A_834 & ~w1374;
assign w13242 = ~A_831 & ~w1379;
assign w13243 = ~A_840 & ~w1422;
assign w13244 = ~A_837 & ~w1427;
assign w13245 = ~A_846 & ~w1456;
assign w13246 = ~A_843 & ~w1461;
assign w13247 = ~A_474 & ~w1589;
assign w13248 = ~A_471 & ~w1591;
assign w13249 = ~A_468 & ~w1622;
assign w13250 = ~A_465 & ~w1624;
assign w13251 = ~A_486 & ~w1658;
assign w13252 = ~A_483 & ~w1660;
assign w13253 = ~A_480 & ~w1691;
assign w13254 = ~A_477 & ~w1693;
assign w13255 = ~A_510 & ~w1730;
assign w13256 = ~A_507 & ~w1732;
assign w13257 = ~A_504 & ~w1763;
assign w13258 = ~A_501 & ~w1765;
assign w13259 = ~A_498 & ~w1799;
assign w13260 = ~A_495 & ~w1801;
assign w13261 = ~A_492 & ~w1832;
assign w13262 = ~A_489 & ~w1834;
assign w13263 = ~A_558 & ~w1874;
assign w13264 = ~A_555 & ~w1876;
assign w13265 = ~A_552 & ~w1907;
assign w13266 = ~A_549 & ~w1909;
assign w13267 = ~A_546 & ~w1943;
assign w13268 = ~A_543 & ~w1945;
assign w13269 = ~A_540 & ~w1976;
assign w13270 = ~A_537 & ~w1978;
assign w13271 = ~A_534 & ~w2015;
assign w13272 = ~A_531 & ~w2017;
assign w13273 = ~A_528 & ~w2048;
assign w13274 = ~A_525 & ~w2050;
assign w13275 = ~A_522 & ~w2084;
assign w13276 = ~A_519 & ~w2086;
assign w13277 = ~A_516 & ~w2117;
assign w13278 = ~A_513 & ~w2119;
assign w13279 = ~A_654 & ~w2162;
assign w13280 = ~A_651 & ~w2164;
assign w13281 = ~A_648 & ~w2195;
assign w13282 = ~A_645 & ~w2197;
assign w13283 = ~A_642 & ~w2231;
assign w13284 = ~A_639 & ~w2233;
assign w13285 = ~A_636 & ~w2264;
assign w13286 = ~A_633 & ~w2266;
assign w13287 = ~A_630 & ~w2303;
assign w13288 = ~A_627 & ~w2305;
assign w13289 = ~A_624 & ~w2336;
assign w13290 = ~A_621 & ~w2338;
assign w13291 = ~A_618 & ~w2372;
assign w13292 = ~A_615 & ~w2374;
assign w13293 = ~A_612 & ~w2405;
assign w13294 = ~A_609 & ~w2407;
assign w13295 = ~A_606 & ~w2447;
assign w13296 = ~A_603 & ~w2449;
assign w13297 = ~A_600 & ~w2480;
assign w13298 = ~A_597 & ~w2482;
assign w13299 = ~A_594 & ~w2516;
assign w13300 = ~A_591 & ~w2518;
assign w13301 = ~A_588 & ~w2549;
assign w13302 = ~A_585 & ~w2551;
assign w13303 = ~A_582 & ~w2588;
assign w13304 = ~A_579 & ~w2590;
assign w13305 = ~A_576 & ~w2621;
assign w13306 = ~A_573 & ~w2623;
assign w13307 = ~A_570 & ~w2657;
assign w13308 = ~A_567 & ~w2659;
assign w13309 = ~A_564 & ~w2690;
assign w13310 = ~A_561 & ~w2692;
assign w13311 = ~A_990 & ~w3279;
assign w13312 = ~A_987 & ~w3284;
assign w13313 = ~A_966 & ~w3364;
assign w13314 = ~A_963 & ~w3366;
assign w13315 = w3622 & w3575;
assign w13316 = w3701 & w3716;
assign w13317 = w3701 & ~w3716;
assign w13318 = w3774 & w3766;
assign w13319 = ~A_5 & ~w3804;
assign w13320 = ~A_2 & ~w3806;
assign w13321 = w3803 & ~w3810;
assign w13322 = w3998 & ~w3919;
assign w13323 = w3919 & ~w3998;
assign w13324 = w4017 & w4003;
assign w13325 = w3919 & w3998;
assign w13326 = w4105 & w4058;
assign w13327 = w4184 & ~w4199;
assign w13328 = w4215 & ~w4025;
assign w13329 = ~w4025 & ~w4231;
assign w13330 = w4218 & w4231;
assign w13331 = ~w4025 & w4231;
assign w13332 = w4218 & ~w4231;
assign w13333 = ~A_942 & ~w4280;
assign w13334 = ~A_939 & ~w4282;
assign w13335 = ~A_936 & ~w4313;
assign w13336 = ~A_933 & ~w4315;
assign w13337 = ~A_930 & ~w4349;
assign w13338 = ~A_927 & ~w4351;
assign w13339 = ~A_924 & ~w4382;
assign w13340 = ~A_921 & ~w4384;
assign w13341 = ~A_918 & ~w4421;
assign w13342 = ~A_915 & ~w4423;
assign w13343 = ~A_912 & ~w4454;
assign w13344 = ~A_909 & ~w4456;
assign w13345 = ~A_906 & ~w4490;
assign w13346 = ~A_903 & ~w4492;
assign w13347 = ~A_900 & ~w4523;
assign w13348 = ~A_897 & ~w4525;
assign w13349 = ~A_894 & ~w4565;
assign w13350 = ~A_891 & ~w4567;
assign w13351 = ~A_888 & ~w4598;
assign w13352 = ~A_885 & ~w4600;
assign w13353 = ~A_882 & ~w4634;
assign w13354 = ~A_879 & ~w4636;
assign w13355 = ~A_876 & ~w4667;
assign w13356 = ~A_873 & ~w4669;
assign w13357 = ~A_870 & ~w4706;
assign w13358 = ~A_867 & ~w4708;
assign w13359 = ~A_864 & ~w4739;
assign w13360 = ~A_861 & ~w4741;
assign w13361 = ~A_858 & ~w4775;
assign w13362 = ~A_855 & ~w4777;
assign w13363 = ~A_852 & ~w4808;
assign w13364 = ~A_849 & ~w4810;
assign w13365 = w5136 & w5089;
assign w13366 = w5215 & ~w5230;
assign w13367 = w5404 & ~w5399;
assign w13368 = w5399 & ~w5404;
assign w13369 = w5423 & w5409;
assign w13370 = w5399 & w5404;
assign w13371 = w5593 & ~w5514;
assign w13372 = w5514 & ~w5593;
assign w13373 = w5612 & w5598;
assign w13374 = w5514 & w5593;
assign w13375 = w5700 & w5653;
assign w13376 = w5779 & ~w5794;
assign w13377 = w5810 & ~w5620;
assign w13378 = ~w5620 & ~w5825;
assign w13379 = w5813 & w5825;
assign w13380 = ~w5620 & w5825;
assign w13381 = w5813 & ~w5825;
assign w13382 = w6434 & ~w6429;
assign w13383 = w6429 & ~w6434;
assign w13384 = w6453 & w6439;
assign w13385 = w6429 & w6434;
assign w13386 = w6477 & w6463;
assign w13387 = w6492 & ~w6497;
assign w13388 = w6512 & w6461;
assign w13389 = w6536 & w6522;
assign w13390 = w6551 & ~w6556;
assign w13391 = w6586 & ~w6581;
assign w13392 = w6581 & ~w6586;
assign w13393 = w6605 & w6591;
assign w13394 = w6581 & w6586;
assign w13395 = w6788 & ~w6709;
assign w13396 = w6709 & ~w6788;
assign w13397 = w6807 & w6793;
assign w13398 = w6709 & w6788;
assign w13399 = w6895 & w6848;
assign w13400 = w6974 & ~w6989;
assign w13401 = w7005 & ~w6815;
assign w13402 = ~w6815 & w7302;
assign w13403 = w7008 & ~w7302;
assign w13404 = w7322 & w7308;
assign w13405 = w7337 & ~w7342;
assign w13406 = w7372 & ~w7367;
assign w13407 = w7367 & ~w7372;
assign w13408 = w7391 & w7377;
assign w13409 = w7367 & w7372;
assign w13410 = ~w6815 & ~w7302;
assign w13411 = w7008 & w7302;
assign w13412 = w7492 & w7445;
assign w13413 = w7571 & ~w7586;
assign w13414 = w7760 & ~w7755;
assign w13415 = w7755 & ~w7760;
assign w13416 = w7779 & w7765;
assign w13417 = w7755 & w7760;
assign w13418 = w7740 & w7787;
assign w13419 = w7968 & w7954;
assign w13420 = w7870 & w7949;
assign w13421 = w8170 & w7975;
assign w13422 = ~w7793 & ~w8197;
assign w13423 = w8199 & ~w7412;
assign w13424 = ~w7412 & ~w8214;
assign w13425 = w8202 & w8214;
assign w13426 = ~w7412 & w8214;
assign w13427 = w8202 & ~w8214;
assign w13428 = w8668 & ~w8258;
assign w13429 = ~w8668 & w8258;
assign w13430 = w3700 & w8304;
assign w13431 = w3622 & w8290;
assign w13432 = w11413 & ~w11415;
assign w13433 = w11417 & ~w11418;
assign w13434 = w11420 & ~w11422;
assign w13435 = w11424 & ~w11426;
assign w13436 = w11428 & ~w11429;
assign w13437 = w10688 & ~w10689;
assign w13438 = w11445 & ~w11448;
assign w13439 = w11450 & ~w11452;
assign w13440 = w11454 & ~w11455;
assign w13441 = w11547 & ~w11548;
assign w13442 = w11550 & ~w11551;
assign w13443 = w11553 & ~w11554;
assign w13444 = w11556 & ~w11559;
assign w13445 = w11561 & ~w11563;
assign w13446 = w11565 & ~w11566;
assign w13447 = w11575 & ~w11578;
assign w13448 = w11580 & ~w11582;
assign w13449 = w11584 & ~w11585;
assign w13450 = w11600 & ~w11601;
assign w13451 = w11603 & ~w11606;
assign w13452 = w11608 & ~w11610;
assign w13453 = w11612 & ~w11613;
assign w13454 = w11622 & ~w11625;
assign w13455 = w11627 & ~w11629;
assign w13456 = w11631 & ~w11632;
assign w13457 = w11653 & ~w11654;
assign w13458 = w11656 & ~w11657;
assign w13459 = w11659 & ~w11662;
assign w13460 = w11664 & ~w11666;
assign w13461 = w11668 & ~w11669;
assign w13462 = w11678 & ~w11681;
assign w13463 = w11683 & ~w11685;
assign w13464 = w11687 & ~w11688;
assign w13465 = w11703 & ~w11704;
assign w13466 = w11706 & ~w11709;
assign w13467 = w11711 & ~w11713;
assign w13468 = w11715 & ~w11716;
assign w13469 = ~w11739 & ~w11721;
assign w13470 = ~w11693 & ~w11674;
assign w13471 = ~w11637 & ~w11618;
assign w13472 = ~w11590 & ~w11571;
assign w13473 = ~w11460 & ~w11441;
assign w13474 = ~w12586 & w8254;
assign w13475 = w12595 & ~w12623;
assign w13476 = w12675 & w12955;
assign w13477 = w12675 & ~w13174;
assign w13478 = w339 & w296;
assign w13479 = ~w355 & ~w340;
assign w13480 = w340 & w355;
assign w13481 = w355 & ~w340;
assign w13482 = w360 & w263;
assign w13483 = w702 & w692;
assign w13484 = ~w708 & ~w703;
assign w13485 = w708 & ~w703;
assign w13486 = w713 & w690;
assign w13487 = w935 & w892;
assign w13488 = ~w951 & ~w936;
assign w13489 = w951 & ~w936;
assign w13490 = w956 & w859;
assign w13491 = w1497 & w1454;
assign w13492 = ~w1513 & ~w1498;
assign w13493 = w1498 & w1513;
assign w13494 = w1513 & ~w1498;
assign w13495 = w1518 & w1421;
assign w13496 = w2758 & w2748;
assign w13497 = ~w2764 & ~w2759;
assign w13498 = w2764 & ~w2759;
assign w13499 = w2769 & w2746;
assign w13500 = w2900 & w2890;
assign w13501 = ~w2906 & ~w2901;
assign w13502 = w2901 & w2906;
assign w13503 = w2906 & ~w2901;
assign w13504 = w2911 & w2888;
assign w13505 = w3015 & w3005;
assign w13506 = ~w3021 & ~w3016;
assign w13507 = w3016 & w3021;
assign w13508 = w3021 & ~w3016;
assign w13509 = w3026 & w3003;
assign w13510 = w3074 & w3064;
assign w13511 = ~w3080 & ~w3075;
assign w13512 = w3080 & ~w3075;
assign w13513 = w3085 & w3062;
assign w13514 = ~A_972 & ~w3163;
assign w13515 = ~A_969 & ~w3168;
assign w13516 = ~A_978 & ~w3197;
assign w13517 = ~A_975 & ~w3202;
assign w13518 = ~A_984 & ~w3245;
assign w13519 = ~A_981 & ~w3250;
assign w13520 = w3320 & w3277;
assign w13521 = w3336 & ~w3321;
assign w13522 = w3341 & w3244;
assign w13523 = ~A_960 & ~w3397;
assign w13524 = ~A_957 & ~w3399;
assign w13525 = ~A_954 & ~w3433;
assign w13526 = ~A_951 & ~w3435;
assign w13527 = ~A_948 & ~w3466;
assign w13528 = ~A_945 & ~w3468;
assign w13529 = w4915 & w4905;
assign w13530 = ~w4921 & ~w4916;
assign w13531 = w4916 & w4921;
assign w13532 = w4921 & ~w4916;
assign w13533 = w4926 & w4903;
assign w13534 = w4974 & w4964;
assign w13535 = ~w4980 & ~w4975;
assign w13536 = w4980 & ~w4975;
assign w13537 = w4985 & w4962;
assign w13538 = w7790 & ~w7787;
assign w13539 = w8262 & ~w8491;
assign w13540 = ~w8493 & w8260;
assign w13541 = w8493 & ~w8260;
assign w13542 = w5020 & w5015;
assign w13543 = w4999 & w4994;
assign w13544 = w4951 & w4946;
assign w13545 = w4969 & w4964;
assign w13546 = w4869 & w4864;
assign w13547 = w4848 & w4843;
assign w13548 = w4892 & w4887;
assign w13549 = w4910 & w4905;
assign w13550 = w3120 & w3115;
assign w13551 = w3099 & w3094;
assign w13552 = w3051 & w3046;
assign w13553 = w3069 & w3064;
assign w13554 = w2969 & w2964;
assign w13555 = w2948 & w2943;
assign w13556 = w2992 & w2987;
assign w13557 = w3010 & w3005;
assign w13558 = w2804 & w2799;
assign w13559 = w2783 & w2778;
assign w13560 = w2735 & w2730;
assign w13561 = w2753 & w2748;
assign w13562 = w2854 & w2849;
assign w13563 = w2833 & w2828;
assign w13564 = w2877 & w2872;
assign w13565 = w2895 & w2890;
assign w13566 = w748 & w743;
assign w13567 = w727 & w722;
assign w13568 = w679 & w674;
assign w13569 = w697 & w692;
assign w13570 = w165 & w160;
assign w13571 = w70 & w32;
assign w13572 = w252 & w214;
assign w13573 = w334 & w296;
assign w13574 = w1135 & w1130;
assign w13575 = w1114 & w1109;
assign w13576 = w848 & w810;
assign w13577 = w930 & w892;
assign w13578 = w1323 & w1318;
assign w13579 = w1228 & w1190;
assign w13580 = w1410 & w1372;
assign w13581 = w1492 & w1454;
assign w13582 = ~w8644 & ~w8630;
assign w13583 = w4883 & ~w10792;
assign w13584 = ~w8608 & ~w8594;
assign w13585 = ~w8564 & ~w8550;
assign w13586 = w5034 & ~w10847;
assign w13587 = ~w8528 & ~w8514;
assign w13588 = ~w10037 & ~w10023;
assign w13589 = w1337 & ~w10934;
assign w13590 = ~w10001 & ~w9987;
assign w13591 = ~w9957 & ~w9943;
assign w13592 = w1149 & ~w10990;
assign w13593 = ~w9921 & ~w9907;
assign w13594 = ~w9869 & ~w9855;
assign w13595 = w179 & ~w11056;
assign w13596 = ~w9833 & ~w9819;
assign w13597 = ~w9789 & ~w9775;
assign w13598 = w762 & ~w11112;
assign w13599 = ~w9753 & ~w9739;
assign w13600 = ~w9693 & ~w9679;
assign w13601 = w2868 & ~w11188;
assign w13602 = ~w9657 & ~w9643;
assign w13603 = ~w9613 & ~w9599;
assign w13604 = w2818 & ~w11244;
assign w13605 = ~w9577 & ~w9563;
assign w13606 = ~w9525 & ~w9511;
assign w13607 = w2983 & ~w11310;
assign w13608 = ~w9489 & ~w9475;
assign w13609 = ~w9445 & ~w9431;
assign w13610 = w3134 & ~w11366;
assign w13611 = ~w9409 & ~w9395;
assign w13612 = ~w12004 & w12002;
assign w13613 = (~w12004 & ~w11728) | (~w12004 & w13612) | (~w11728 & w13612);
assign w13614 = ~w12009 & w12008;
assign w13615 = (~w12009 & ~w11709) | (~w12009 & w13614) | (~w11709 & w13614);
assign w13616 = ~w12027 & w12025;
assign w13617 = (~w12027 & ~w11681) | (~w12027 & w13616) | (~w11681 & w13616);
assign w13618 = ~w12032 & w12031;
assign w13619 = (~w12032 & ~w11662) | (~w12032 & w13618) | (~w11662 & w13618);
assign w13620 = ~w12059 & w12057;
assign w13621 = (~w12059 & ~w11625) | (~w12059 & w13620) | (~w11625 & w13620);
assign w13622 = ~w12064 & w12063;
assign w13623 = (~w12064 & ~w11606) | (~w12064 & w13622) | (~w11606 & w13622);
assign w13624 = ~w12082 & w12080;
assign w13625 = (~w12082 & ~w11578) | (~w12082 & w13624) | (~w11578 & w13624);
assign w13626 = ~w12087 & w12086;
assign w13627 = (~w12087 & ~w11559) | (~w12087 & w13626) | (~w11559 & w13626);
assign w13628 = ~w12126 & w12124;
assign w13629 = (~w12126 & ~w11448) | (~w12126 & w13628) | (~w11448 & w13628);
assign w13630 = ~w11439 & w11437;
assign w13631 = (~w11439 & ~w10689) | (~w11439 & w13630) | (~w10689 & w13630);
assign w13632 = ~w12133 & w12139;
assign w13633 = w12146 & ~w12143;
assign w13634 = w12300 & ~w12302;
assign w13635 = w12304 & ~w12305;
assign w13636 = w12307 & ~w12309;
assign w13637 = w12316 & ~w12318;
assign w13638 = w12335 & ~w12336;
assign w13639 = w12338 & ~w12341;
assign w13640 = w12345 & ~w12347;
assign w13641 = w12351 & ~w12352;
assign w13642 = w12361 & ~w12364;
assign w13643 = w12368 & ~w12370;
assign w13644 = w12374 & ~w12375;
assign w13645 = ~w12380 & ~w12357;
assign w13646 = w12682 & w12684;
assign w13647 = (w12680 & w14049) | (w12680 & w14050) | (w14049 & w14050);
assign w13648 = w12688 & w12692;
assign w13649 = w12693 & w12701;
assign w13650 = w12679 & w12963;
assign w13651 = ~w12643 & w12689;
assign w13652 = ~w12643 & ~w12965;
assign w13653 = w75 & w32;
assign w13654 = w155 & ~w76;
assign w13655 = w76 & ~w155;
assign w13656 = ~w155 & ~w76;
assign w13657 = w178 & ~w176;
assign w13658 = w261 & w214;
assign w13659 = w340 & ~w355;
assign w13660 = w376 & w181;
assign w13661 = w688 & w674;
assign w13662 = w703 & w708;
assign w13663 = w703 & ~w708;
assign w13664 = w732 & w722;
assign w13665 = w738 & ~w733;
assign w13666 = w733 & ~w738;
assign w13667 = ~w738 & ~w733;
assign w13668 = w761 & ~w759;
assign w13669 = w857 & w810;
assign w13670 = w936 & w951;
assign w13671 = w936 & ~w951;
assign w13672 = w1119 & w1109;
assign w13673 = w1125 & ~w1120;
assign w13674 = w1120 & ~w1125;
assign w13675 = ~w1125 & ~w1120;
assign w13676 = w1148 & ~w1146;
assign w13677 = w1233 & w1190;
assign w13678 = w1313 & ~w1234;
assign w13679 = w1234 & ~w1313;
assign w13680 = ~w1313 & ~w1234;
assign w13681 = w1336 & ~w1334;
assign w13682 = w1419 & w1372;
assign w13683 = w1498 & ~w1513;
assign w13684 = w1529 & ~w1339;
assign w13685 = ~w1339 & ~w1544;
assign w13686 = w1532 & w1544;
assign w13687 = ~w1339 & w1544;
assign w13688 = w1532 & ~w1544;
assign w13689 = w2744 & w2730;
assign w13690 = w2759 & w2764;
assign w13691 = w2759 & ~w2764;
assign w13692 = w2788 & w2778;
assign w13693 = w2794 & ~w2789;
assign w13694 = w2789 & ~w2794;
assign w13695 = ~w2794 & ~w2789;
assign w13696 = w2817 & ~w2815;
assign w13697 = w2838 & w2828;
assign w13698 = w2844 & ~w2839;
assign w13699 = w2839 & ~w2844;
assign w13700 = ~w2844 & ~w2839;
assign w13701 = w2867 & ~w2865;
assign w13702 = w2886 & w2872;
assign w13703 = w2901 & ~w2906;
assign w13704 = w2916 & ~w2870;
assign w13705 = ~w2870 & ~w2925;
assign w13706 = ~w2870 & w2925;
assign w13707 = w2919 & ~w2925;
assign w13708 = w2953 & w2943;
assign w13709 = w2959 & ~w2954;
assign w13710 = w2954 & ~w2959;
assign w13711 = ~w2959 & ~w2954;
assign w13712 = w2982 & ~w2980;
assign w13713 = w3001 & w2987;
assign w13714 = w3016 & ~w3021;
assign w13715 = w3036 & w2985;
assign w13716 = w3060 & w3046;
assign w13717 = w3075 & w3080;
assign w13718 = w3075 & ~w3080;
assign w13719 = w3104 & w3094;
assign w13720 = w3110 & ~w3105;
assign w13721 = w3105 & ~w3110;
assign w13722 = ~w3110 & ~w3105;
assign w13723 = w3133 & ~w3131;
assign w13724 = w3242 & w3195;
assign w13725 = ~w3336 & ~w3321;
assign w13726 = w3321 & w3336;
assign w13727 = w3321 & ~w3336;
assign w13728 = w3504 & w3494;
assign w13729 = w3510 & ~w3505;
assign w13730 = w3505 & ~w3510;
assign w13731 = ~w3510 & ~w3505;
assign w13732 = w3533 & ~w3531;
assign w13733 = w3520 & w3515;
assign w13734 = w3499 & w3494;
assign w13735 = w3233 & w3195;
assign w13736 = w3315 & w3277;
assign w13737 = w10911 & ~w10914;
assign w13738 = w1497 & w10031;
assign w13739 = w1419 & w10017;
assign w13740 = w1233 & w9995;
assign w13741 = w1332 & w9981;
assign w13742 = w10967 & ~w10970;
assign w13743 = w935 & w9951;
assign w13744 = w857 & w9937;
assign w13745 = w1119 & w9915;
assign w13746 = w1144 & w9901;
assign w13747 = w11033 & ~w11036;
assign w13748 = w339 & w9863;
assign w13749 = w261 & w9849;
assign w13750 = w75 & w9827;
assign w13751 = w174 & w9813;
assign w13752 = w11089 & ~w11092;
assign w13753 = w702 & w9783;
assign w13754 = w688 & w9769;
assign w13755 = w732 & w9747;
assign w13756 = w757 & w9733;
assign w13757 = w11165 & ~w11168;
assign w13758 = w2900 & w9687;
assign w13759 = w2886 & w9673;
assign w13760 = w2838 & w9651;
assign w13761 = w2863 & w9637;
assign w13762 = w11221 & ~w11224;
assign w13763 = w2758 & w9607;
assign w13764 = w2744 & w9593;
assign w13765 = w2788 & w9571;
assign w13766 = w2813 & w9557;
assign w13767 = w11287 & ~w11290;
assign w13768 = w3015 & w9519;
assign w13769 = w3001 & w9505;
assign w13770 = w2953 & w9483;
assign w13771 = w2978 & w9469;
assign w13772 = w11343 & ~w11346;
assign w13773 = w3074 & w9439;
assign w13774 = w3060 & w9425;
assign w13775 = w3104 & w9403;
assign w13776 = w3129 & w9389;
assign w13777 = ~w11384 & ~w11361;
assign w13778 = ~w11328 & ~w11305;
assign w13779 = ~w11262 & ~w11239;
assign w13780 = ~w11206 & ~w11183;
assign w13781 = ~w11130 & ~w11107;
assign w13782 = ~w11074 & ~w11051;
assign w13783 = ~w11008 & ~w10985;
assign w13784 = ~w10952 & ~w10929;
assign w13785 = w11454 & w12122;
assign w13786 = ~w12133 & ~w12139;
assign w13787 = w12316 & w12326;
assign w13788 = w12327 & ~w12315;
assign w13789 = w12449 & ~w12451;
assign w13790 = w12453 & ~w12454;
assign w13791 = w12330 & ~w12328;
assign w13792 = w12330 & w12458;
assign w13793 = w12461 & ~w12464;
assign w13794 = w12468 & ~w12470;
assign w13795 = w12474 & ~w12475;
assign w13796 = ~w12457 & ~w12480;
assign w13797 = w174 & w160;
assign w13798 = w76 & w155;
assign w13799 = w371 & ~w181;
assign w13800 = w757 & w743;
assign w13801 = w733 & w738;
assign w13802 = w718 & w764;
assign w13803 = w767 & ~w764;
assign w13804 = w1144 & w1130;
assign w13805 = w1120 & w1125;
assign w13806 = w1105 & w1151;
assign w13807 = w1154 & ~w1151;
assign w13808 = w1332 & w1318;
assign w13809 = w1234 & w1313;
assign w13810 = w1534 & w1339;
assign w13811 = ~w1157 & ~w1561;
assign w13812 = w1563 & ~w777;
assign w13813 = ~w777 & w2724;
assign w13814 = w1566 & ~w2724;
assign w13815 = w2813 & w2799;
assign w13816 = w2789 & w2794;
assign w13817 = w2774 & w2820;
assign w13818 = w2823 & ~w2820;
assign w13819 = w2863 & w2849;
assign w13820 = w2839 & w2844;
assign w13821 = w2921 & w2870;
assign w13822 = ~w2826 & w2937;
assign w13823 = w2978 & w2964;
assign w13824 = w2954 & w2959;
assign w13825 = w3031 & ~w2985;
assign w13826 = w3129 & w3115;
assign w13827 = w3105 & w3110;
assign w13828 = w3090 & w3136;
assign w13829 = w3139 & ~w3136;
assign w13830 = w2939 & w3149;
assign w13831 = ~w777 & ~w2724;
assign w13832 = w1566 & w2724;
assign w13833 = w3529 & w3515;
assign w13834 = w3505 & w3510;
assign w13835 = w3490 & w3536;
assign w13836 = w3539 & ~w3536;
assign w13837 = ~A_996 & ~w3744;
assign w13838 = ~A_993 & ~w3746;
assign w13839 = ~A_999 & ~w3817;
assign w13840 = w3797 & w3836;
assign w13841 = w3839 & ~w3836;
assign w13842 = w4220 & w4025;
assign w13843 = ~w3842 & ~w4248;
assign w13844 = w4250 & ~w3542;
assign w13845 = ~w3842 & w4248;
assign w13846 = w4256 & w3542;
assign w13847 = w4853 & w4843;
assign w13848 = w4859 & ~w4854;
assign w13849 = w4854 & ~w4859;
assign w13850 = w4878 & w4864;
assign w13851 = ~w4859 & ~w4854;
assign w13852 = w4882 & ~w4880;
assign w13853 = w4901 & w4887;
assign w13854 = w4916 & ~w4921;
assign w13855 = w4931 & ~w4885;
assign w13856 = ~w4885 & w4940;
assign w13857 = w4934 & ~w4940;
assign w13858 = w4960 & w4946;
assign w13859 = w4975 & w4980;
assign w13860 = w4975 & ~w4980;
assign w13861 = w5004 & w4994;
assign w13862 = w5010 & ~w5005;
assign w13863 = w5005 & ~w5010;
assign w13864 = w5029 & w5015;
assign w13865 = ~w5010 & ~w5005;
assign w13866 = w5033 & ~w5031;
assign w13867 = w4990 & w5036;
assign w13868 = ~w4885 & ~w4940;
assign w13869 = w4934 & w4940;
assign w13870 = w5384 & w5431;
assign w13871 = w5434 & ~w5431;
assign w13872 = w5815 & w5620;
assign w13873 = ~w5437 & w6412;
assign w13874 = w6507 & ~w6461;
assign w13875 = w6566 & w6613;
assign w13876 = w6616 & ~w6613;
assign w13877 = w6414 & w6626;
assign w13878 = w7010 & w6815;
assign w13879 = w7352 & w7399;
assign w13880 = w7402 & ~w7399;
assign w13881 = ~w7793 & w8197;
assign w13882 = w8204 & w7412;
assign w13883 = (~w8232 & w6631) | (~w8232 & w14051) | (w6631 & w14051);
assign w13884 = w8234 & ~w5056;
assign w13885 = (w8232 & w6631) | (w8232 & w14052) | (w6631 & w14052);
assign w13886 = w8246 & w5056;
assign w13887 = w8237 & ~w3162;
assign w13888 = w10071 & ~w8254;
assign w13889 = w8673 & ~w8256;
assign w13890 = w8262 & w8491;
assign w13891 = w8260 & ~w10593;
assign w13892 = (~w8275 & w8268) | (~w8275 & w14053) | (w8268 & w14053);
assign w13893 = ~w10661 & ~w12949;
assign w13894 = ~w8475 & ~w8461;
assign w13895 = w3320 & w8469;
assign w13896 = w3242 & w8455;
assign w13897 = w10707 & ~w10720;
assign w13898 = ~w8439 & ~w8425;
assign w13899 = w3504 & w8433;
assign w13900 = w3529 & w8419;
assign w13901 = w10729 & ~w10742;
assign w13902 = w10769 & ~w10772;
assign w13903 = w4915 & w8638;
assign w13904 = w4901 & w8624;
assign w13905 = w4853 & w8602;
assign w13906 = w4878 & w8588;
assign w13907 = w10821 & ~w10822;
assign w13908 = w10824 & ~w10827;
assign w13909 = w4974 & w8558;
assign w13910 = w4960 & w8544;
assign w13911 = w5004 & w8522;
assign w13912 = w5029 & w8508;
assign w13913 = w10594 & ~w10881;
assign w13914 = w10078 & w11412;
assign w13915 = w10594 & w10881;
assign w13916 = ~w10661 & ~w11435;
assign w13917 = ~w10743 & ~w10721;
assign w13918 = w10707 & ~w11473;
assign w13919 = w10729 & ~w11477;
assign w13920 = w11472 & ~w11482;
assign w13921 = w11494 & ~w11495;
assign w13922 = ~w10865 & ~w10842;
assign w13923 = w11501 & ~w11503;
assign w13924 = w11505 & ~w11506;
assign w13925 = w11500 & ~w11510;
assign w13926 = ~w10810 & ~w10787;
assign w13927 = w11519 & ~w11521;
assign w13928 = w11523 & ~w11524;
assign w13929 = w11518 & ~w11528;
assign w13930 = w11781 & ~w11783;
assign w13931 = w11785 & ~w11786;
assign w13932 = w11800 & ~w11802;
assign w13933 = w11804 & ~w11805;
assign w13934 = w11828 & ~w11830;
assign w13935 = w11832 & ~w11833;
assign w13936 = w11847 & ~w11849;
assign w13937 = w11851 & ~w11852;
assign w13938 = w11884 & ~w11886;
assign w13939 = w11888 & ~w11889;
assign w13940 = w11903 & ~w11905;
assign w13941 = w11907 & ~w11908;
assign w13942 = w11931 & ~w11933;
assign w13943 = w11935 & ~w11936;
assign w13944 = w11950 & ~w11952;
assign w13945 = w11954 & ~w11955;
assign w13946 = w11733 & w12000;
assign w13947 = w11715 & w12006;
assign w13948 = w11687 & w12023;
assign w13949 = w11668 & w12029;
assign w13950 = w11631 & w12055;
assign w13951 = w11612 & w12061;
assign w13952 = w11584 & w12078;
assign w13953 = w11565 & w12084;
assign w13954 = ~w12138 & w12137;
assign w13955 = (~w12138 & ~w11472) | (~w12138 & w13954) | (~w11472 & w13954);
assign w13956 = ~w11529 & ~w11511;
assign w13957 = w11523 & w12154;
assign w13958 = w11518 & ~w12156;
assign w13959 = ~w12158 & w12156;
assign w13960 = (~w12158 & ~w11518) | (~w12158 & w13959) | (~w11518 & w13959);
assign w13961 = w11505 & w12160;
assign w13962 = w11500 & ~w12162;
assign w13963 = ~w12163 & w12162;
assign w13964 = (~w12163 & ~w11500) | (~w12163 & w13963) | (~w11500 & w13963);
assign w13965 = w12185 & ~w12186;
assign w13966 = w12188 & ~w12189;
assign w13967 = ~w11960 & ~w11941;
assign w13968 = w11954 & w12195;
assign w13969 = w12197 & ~w12199;
assign w13970 = w11935 & w12201;
assign w13971 = w12203 & ~w12204;
assign w13972 = w12194 & ~w12208;
assign w13973 = ~w11913 & ~w11894;
assign w13974 = w11907 & w12217;
assign w13975 = w12219 & ~w12221;
assign w13976 = w11888 & w12223;
assign w13977 = w12225 & ~w12226;
assign w13978 = w12216 & ~w12230;
assign w13979 = w12241 & ~w12242;
assign w13980 = ~w11857 & ~w11838;
assign w13981 = w11851 & w12248;
assign w13982 = w12250 & ~w12252;
assign w13983 = w11832 & w12254;
assign w13984 = w12256 & ~w12257;
assign w13985 = w12247 & ~w12261;
assign w13986 = ~w11810 & ~w11791;
assign w13987 = w11804 & w12270;
assign w13988 = w12272 & ~w12274;
assign w13989 = w11785 & w12276;
assign w13990 = w12278 & ~w12279;
assign w13991 = w12269 & ~w12283;
assign w13992 = w12313 & ~w12314;
assign w13993 = w12322 & ~w12323;
assign w13994 = w12396 & ~w12397;
assign w13995 = ~w12284 & ~w12262;
assign w13996 = w12256 & w12403;
assign w13997 = w12247 & ~w12405;
assign w13998 = ~w12407 & w12405;
assign w13999 = (~w12407 & ~w12247) | (~w12407 & w13998) | (~w12247 & w13998);
assign w14000 = w12278 & w12409;
assign w14001 = w12269 & ~w12411;
assign w14002 = ~w12412 & w12411;
assign w14003 = (~w12412 & ~w12269) | (~w12412 & w14002) | (~w12269 & w14002);
assign w14004 = w12402 & ~w12416;
assign w14005 = ~w12231 & ~w12209;
assign w14006 = w12203 & w12425;
assign w14007 = w12194 & ~w12427;
assign w14008 = ~w12429 & w12427;
assign w14009 = (~w12429 & ~w12194) | (~w12429 & w14008) | (~w12194 & w14008);
assign w14010 = w12225 & w12431;
assign w14011 = w12216 & ~w12433;
assign w14012 = ~w12434 & w12433;
assign w14013 = (~w12434 & ~w12216) | (~w12434 & w14012) | (~w12216 & w14012);
assign w14014 = w12424 & ~w12438;
assign w14015 = w12456 & w12328;
assign w14016 = w12456 & ~w13791;
assign w14017 = w12374 & w12466;
assign w14018 = w12351 & w12472;
assign w14019 = ~w12439 & ~w12417;
assign w14020 = w12424 & ~w12497;
assign w14021 = ~w12499 & w12497;
assign w14022 = (~w12499 & ~w12424) | (~w12499 & w14021) | (~w12424 & w14021);
assign w14023 = w12402 & ~w12503;
assign w14024 = ~w12504 & w12503;
assign w14025 = (~w12504 & ~w12402) | (~w12504 & w14024) | (~w12402 & w14024);
assign w14026 = w12494 & ~w12508;
assign w14027 = w12513 & ~w12516;
assign w14028 = w12484 & ~w12486;
assign w14029 = w12474 & w12520;
assign w14030 = w12522 & ~w12524;
assign w14031 = ~w12537 & w12536;
assign w14032 = (~w12537 & ~w12494) | (~w12537 & w14031) | (~w12494 & w14031);
assign w14033 = ~w12531 & ~w12538;
assign w14034 = w12539 & ~w12541;
assign w14035 = w12526 & ~w12528;
assign w14036 = w12539 & w12545;
assign w14037 = ~w12531 & w12538;
assign w14038 = w12551 & ~w12548;
assign w14039 = w10078 & ~w11412;
assign w14040 = w12586 & ~w8254;
assign w14041 = w8254 & w12593;
assign w14042 = (w12593 & w14041) | (w12593 & ~w12586) | (w14041 & ~w12586);
assign w14043 = ~w3162 & w12593;
assign w14044 = w12615 & ~w12542;
assign w14045 = w8242 & A_1000;
assign w14046 = ~w12646 & ~w12614;
assign w14047 = w12627 & w12664;
assign w14048 = w12684 & w14054;
assign w14049 = w12687 & w12684;
assign w14050 = w12687 & w13646;
assign w14051 = w6627 & ~w8232;
assign w14052 = w6627 & w8232;
assign w14053 = w8270 & ~w8275;
assign w14054 = w12690 & w12682;
assign w14055 = ~w1157 & w1561;
assign w14056 = w1568 & w777;
assign w14057 = ~w2826 & ~w2937;
assign w14058 = w3152 & ~w3149;
assign w14059 = w4854 & w4859;
assign w14060 = w4936 & w4885;
assign w14061 = w5005 & w5010;
assign w14062 = w5039 & ~w5036;
assign w14063 = ~w5437 & ~w6412;
assign w14064 = w6629 & ~w6626;
assign w14065 = w8256 & w10071;
assign w14066 = ~w12614 & w14048;
assign w14067 = ~w12614 & w12964;
assign w14068 = (w11477 & ~w13919) | (w11477 & ~w10727) | (~w13919 & ~w10727);
assign w14069 = (w12162 & ~w13962) | (w12162 & ~w11498) | (~w13962 & ~w11498);
assign w14070 = (w11437 & ~w13168) | (w11437 & ~w11431) | (~w13168 & ~w11431);
assign w14071 = (w12063 & ~w13160) | (w12063 & ~w11604) | (~w13160 & ~w11604);
assign w14072 = (w12086 & ~w13163) | (w12086 & ~w11557) | (~w13163 & ~w11557);
assign w14073 = (w12008 & ~w13153) | (w12008 & ~w11707) | (~w13153 & ~w11707);
assign w14074 = (w12031 & ~w13156) | (w12031 & ~w11660) | (~w13156 & ~w11660);
assign w14075 = (w12433 & ~w14011) | (w12433 & ~w12214) | (~w14011 & ~w12214);
assign w14076 = (w12411 & ~w14001) | (w12411 & ~w12267) | (~w14001 & ~w12267);
assign w14077 = (w12503 & ~w14023) | (w12503 & ~w12400) | (~w14023 & ~w12400);
assign one = 1;
assign maj = ~w12703;// level 60
endmodule

// Benchmark "i5" written by ABC on Sun Apr 22 21:43:04 2018

module i5 ( 
    pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008, pi009,
    pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018, pi019,
    pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028, pi029,
    pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038, pi039,
    pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048, pi049,
    pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058, pi059,
    pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068, pi069,
    pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078, pi079,
    pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088, pi089,
    pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098, pi099,
    pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109,
    pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118, pi119,
    pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128, pi129,
    pi130, pi131, pi132,
    po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10, po11,
    po12, po13, po14, po15, po16, po17, po18, po19, po20, po21, po22, po23,
    po24, po25, po26, po27, po28, po29, po30, po31, po32, po33, po34, po35,
    po36, po37, po38, po39, po40, po41, po42, po43, po44, po45, po46, po47,
    po48, po49, po50, po51, po52, po53, po54, po55, po56, po57, po58, po59,
    po60, po61, po62, po63, po64, po65  );
  input  pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008,
    pi009, pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018,
    pi019, pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028,
    pi029, pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038,
    pi039, pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048,
    pi049, pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058,
    pi059, pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068,
    pi069, pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078,
    pi079, pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088,
    pi089, pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098,
    pi099, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108,
    pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118,
    pi119, pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128,
    pi129, pi130, pi131, pi132;
  output po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10,
    po11, po12, po13, po14, po15, po16, po17, po18, po19, po20, po21, po22,
    po23, po24, po25, po26, po27, po28, po29, po30, po31, po32, po33, po34,
    po35, po36, po37, po38, po39, po40, po41, po42, po43, po44, po45, po46,
    po47, po48, po49, po50, po51, po52, po53, po54, po55, po56, po57, po58,
    po59, po60, po61, po62, po63, po64, po65;
  wire n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
    n211, n212, n214, n215, n216, n217, n219, n221, n222, n223, n224, n225,
    n226, n228, n229, n230, n231, n232, n233, n234, n235, n237, n238, n239,
    n240, n241, n242, n243, n244, n246, n247, n249, n251, n252, n254, n255,
    n256, n257, n258, n259, n260, n261, n263, n264, n266, n268, n270, n271,
    n272, n273, n274, n275, n276, n277, n279, n280, n282, n284, n285, n286,
    n287, n288, n289, n290, n291, n293, n294, n296, n298, n299, n301, n302,
    n303, n304, n305, n306, n307, n308, n310, n311, n312, n313, n314, n315,
    n316, n317, n319, n320, n322, n324, n325, n327, n328, n329, n330, n331,
    n332, n333, n334, n336, n337, n339, n341, n343, n344, n345, n346, n347,
    n348, n349, n350, n352, n353, n355, n357, n358, n359, n360, n361, n362,
    n363, n364, n366, n367, n369, n371, n373, n374, n375, n376, n377, n378,
    n379, n380, n382, n383, n384, n385, n386, n387, n388, n389, n391, n392,
    n394, n396, n397, n399, n400, n401, n402, n403, n404, n405, n406, n408,
    n409, n411, n413, n415, n416, n417, n418, n419, n420, n421, n422, n424,
    n425, n427, n429, n430, n431, n432, n433, n434, n435, n436, n438, n439,
    n441, n443, n444, n445, n446, n447, n448, n449, n450, n452, n453, n454,
    n455, n456, n457, n458, n459, n461, n462, n464, n466, n467, n469, n470,
    n471, n472, n473, n474, n475, n476, n478, n479, n481, n483, n485, n486,
    n487, n488, n489, n490, n491, n492, n494, n495, n497, n499, n500, n501,
    n502, n503, n504, n505, n506, n508, n509, n511;
  assign n200 = pi095 & pi129;
  assign n201 = pi125 & n200;
  assign n202 = pi127 & n201;
  assign n203 = pi131 & n202;
  assign n204 = pi127 & pi128;
  assign n205 = pi125 & n204;
  assign n206 = pi125 & pi126;
  assign n207 = pi125 & pi129;
  assign n208 = pi130 & n207;
  assign n209 = pi127 & n208;
  assign n210 = ~n203 & ~n205;
  assign n211 = ~pi132 & n210;
  assign n212 = ~n206 & ~n209;
  assign po62 = ~n211 | ~n212;
  assign n214 = pi000 & po62;
  assign n215 = pi002 & n214;
  assign n216 = pi000 & pi001;
  assign n217 = ~pi003 & ~n215;
  assign po00 = n216 | ~n217;
  assign n219 = pi002 & po62;
  assign po01 = pi001 | n219;
  assign n221 = pi127 & n200;
  assign n222 = pi131 & n221;
  assign n223 = pi129 & pi130;
  assign n224 = pi127 & n223;
  assign n225 = ~n204 & ~n222;
  assign n226 = ~pi126 & ~n224;
  assign po63 = ~n225 | ~n226;
  assign n228 = pi103 & po63;
  assign n229 = pi101 & n228;
  assign n230 = pi105 & n229;
  assign n231 = pi101 & pi102;
  assign n232 = pi103 & pi104;
  assign n233 = pi101 & n232;
  assign n234 = ~n230 & ~n231;
  assign n235 = ~pi121 & ~n233;
  assign po50 = ~n234 | ~n235;
  assign n237 = pi006 & po50;
  assign n238 = pi004 & n237;
  assign n239 = pi008 & n238;
  assign n240 = pi004 & pi005;
  assign n241 = pi006 & pi007;
  assign n242 = pi004 & n241;
  assign n243 = ~n239 & ~n240;
  assign n244 = ~pi024 & ~n242;
  assign po02 = ~n243 | ~n244;
  assign n246 = pi008 & n237;
  assign n247 = ~pi005 & ~n246;
  assign po03 = n241 | ~n247;
  assign n249 = pi008 & po50;
  assign po04 = pi007 | n249;
  assign n251 = pi105 & n228;
  assign n252 = ~pi102 & ~n251;
  assign po51 = n232 | ~n252;
  assign n254 = pi011 & po51;
  assign n255 = pi009 & n254;
  assign n256 = pi013 & n255;
  assign n257 = pi009 & pi010;
  assign n258 = pi011 & pi012;
  assign n259 = pi009 & n258;
  assign n260 = ~n256 & ~n257;
  assign n261 = ~pi025 & ~n259;
  assign po05 = ~n260 | ~n261;
  assign n263 = pi013 & n254;
  assign n264 = ~pi010 & ~n263;
  assign po06 = n258 | ~n264;
  assign n266 = pi013 & po51;
  assign po07 = pi012 | n266;
  assign n268 = pi105 & po63;
  assign po52 = pi104 | n268;
  assign n270 = pi016 & po52;
  assign n271 = pi014 & n270;
  assign n272 = pi018 & n271;
  assign n273 = pi014 & pi015;
  assign n274 = pi016 & pi017;
  assign n275 = pi014 & n274;
  assign n276 = ~n272 & ~n273;
  assign n277 = ~pi026 & ~n275;
  assign po08 = ~n276 | ~n277;
  assign n279 = pi018 & n270;
  assign n280 = ~pi015 & ~n279;
  assign po09 = n274 | ~n280;
  assign n282 = pi018 & po52;
  assign po10 = pi017 | n282;
  assign n284 = pi021 & po63;
  assign n285 = pi019 & n284;
  assign n286 = pi023 & n285;
  assign n287 = pi019 & pi020;
  assign n288 = pi021 & pi022;
  assign n289 = pi019 & n288;
  assign n290 = ~n286 & ~n287;
  assign n291 = ~pi027 & ~n289;
  assign po11 = ~n290 | ~n291;
  assign n293 = pi023 & n284;
  assign n294 = ~pi020 & ~n293;
  assign po12 = n288 | ~n294;
  assign n296 = pi023 & po63;
  assign po13 = pi022 | n296;
  assign n298 = pi131 & n200;
  assign n299 = ~pi128 & ~n298;
  assign po64 = n223 | ~n299;
  assign n301 = pi108 & po64;
  assign n302 = pi106 & n301;
  assign n303 = pi110 & n302;
  assign n304 = pi106 & pi107;
  assign n305 = pi108 & pi109;
  assign n306 = pi106 & n305;
  assign n307 = ~n303 & ~n304;
  assign n308 = ~pi122 & ~n306;
  assign po53 = ~n307 | ~n308;
  assign n310 = pi030 & po53;
  assign n311 = pi028 & n310;
  assign n312 = pi032 & n311;
  assign n313 = pi028 & pi029;
  assign n314 = pi030 & pi031;
  assign n315 = pi028 & n314;
  assign n316 = ~n312 & ~n313;
  assign n317 = ~pi048 & ~n315;
  assign po14 = ~n316 | ~n317;
  assign n319 = pi032 & n310;
  assign n320 = ~pi029 & ~n319;
  assign po15 = n314 | ~n320;
  assign n322 = pi032 & po53;
  assign po16 = pi031 | n322;
  assign n324 = pi110 & n301;
  assign n325 = ~pi107 & ~n324;
  assign po54 = n305 | ~n325;
  assign n327 = pi035 & po54;
  assign n328 = pi033 & n327;
  assign n329 = pi037 & n328;
  assign n330 = pi033 & pi034;
  assign n331 = pi035 & pi036;
  assign n332 = pi033 & n331;
  assign n333 = ~n329 & ~n330;
  assign n334 = ~pi049 & ~n332;
  assign po17 = ~n333 | ~n334;
  assign n336 = pi037 & n327;
  assign n337 = ~pi034 & ~n336;
  assign po18 = n331 | ~n337;
  assign n339 = pi037 & po54;
  assign po19 = pi036 | n339;
  assign n341 = pi110 & po64;
  assign po55 = pi109 | n341;
  assign n343 = pi040 & po55;
  assign n344 = pi038 & n343;
  assign n345 = pi042 & n344;
  assign n346 = pi038 & pi039;
  assign n347 = pi040 & pi041;
  assign n348 = pi038 & n347;
  assign n349 = ~n345 & ~n346;
  assign n350 = ~pi050 & ~n348;
  assign po20 = ~n349 | ~n350;
  assign n352 = pi042 & n343;
  assign n353 = ~pi039 & ~n352;
  assign po21 = n347 | ~n353;
  assign n355 = pi042 & po55;
  assign po22 = pi041 | n355;
  assign n357 = pi045 & po64;
  assign n358 = pi043 & n357;
  assign n359 = pi047 & n358;
  assign n360 = pi043 & pi044;
  assign n361 = pi045 & pi046;
  assign n362 = pi043 & n361;
  assign n363 = ~n359 & ~n360;
  assign n364 = ~pi051 & ~n362;
  assign po23 = ~n363 | ~n364;
  assign n366 = pi047 & n357;
  assign n367 = ~pi044 & ~n366;
  assign po24 = n361 | ~n367;
  assign n369 = pi047 & po64;
  assign po25 = pi046 | n369;
  assign n371 = pi095 & pi131;
  assign po65 = pi130 | n371;
  assign n373 = pi113 & po65;
  assign n374 = pi111 & n373;
  assign n375 = pi115 & n374;
  assign n376 = pi111 & pi112;
  assign n377 = pi113 & pi114;
  assign n378 = pi111 & n377;
  assign n379 = ~n375 & ~n376;
  assign n380 = ~pi123 & ~n378;
  assign po56 = ~n379 | ~n380;
  assign n382 = pi054 & po56;
  assign n383 = pi052 & n382;
  assign n384 = pi056 & n383;
  assign n385 = pi052 & pi053;
  assign n386 = pi054 & pi055;
  assign n387 = pi052 & n386;
  assign n388 = ~n384 & ~n385;
  assign n389 = ~pi072 & ~n387;
  assign po26 = ~n388 | ~n389;
  assign n391 = pi056 & n382;
  assign n392 = ~pi053 & ~n391;
  assign po27 = n386 | ~n392;
  assign n394 = pi056 & po56;
  assign po28 = pi055 | n394;
  assign n396 = pi115 & n373;
  assign n397 = ~pi112 & ~n396;
  assign po57 = n377 | ~n397;
  assign n399 = pi059 & po57;
  assign n400 = pi057 & n399;
  assign n401 = pi061 & n400;
  assign n402 = pi057 & pi058;
  assign n403 = pi059 & pi060;
  assign n404 = pi057 & n403;
  assign n405 = ~n401 & ~n402;
  assign n406 = ~pi073 & ~n404;
  assign po29 = ~n405 | ~n406;
  assign n408 = pi061 & n399;
  assign n409 = ~pi058 & ~n408;
  assign po30 = n403 | ~n409;
  assign n411 = pi061 & po57;
  assign po31 = pi060 | n411;
  assign n413 = pi115 & po65;
  assign po58 = pi114 | n413;
  assign n415 = pi064 & po58;
  assign n416 = pi062 & n415;
  assign n417 = pi066 & n416;
  assign n418 = pi062 & pi063;
  assign n419 = pi064 & pi065;
  assign n420 = pi062 & n419;
  assign n421 = ~n417 & ~n418;
  assign n422 = ~pi074 & ~n420;
  assign po32 = ~n421 | ~n422;
  assign n424 = pi066 & n415;
  assign n425 = ~pi063 & ~n424;
  assign po33 = n419 | ~n425;
  assign n427 = pi066 & po58;
  assign po34 = pi065 | n427;
  assign n429 = pi069 & po65;
  assign n430 = pi067 & n429;
  assign n431 = pi071 & n430;
  assign n432 = pi067 & pi068;
  assign n433 = pi069 & pi070;
  assign n434 = pi067 & n433;
  assign n435 = ~n431 & ~n432;
  assign n436 = ~pi075 & ~n434;
  assign po35 = ~n435 | ~n436;
  assign n438 = pi071 & n429;
  assign n439 = ~pi068 & ~n438;
  assign po36 = n433 | ~n439;
  assign n441 = pi071 & po65;
  assign po37 = pi070 | n441;
  assign n443 = pi095 & pi118;
  assign n444 = pi116 & n443;
  assign n445 = pi120 & n444;
  assign n446 = pi116 & pi117;
  assign n447 = pi118 & pi119;
  assign n448 = pi116 & n447;
  assign n449 = ~n445 & ~n446;
  assign n450 = ~pi124 & ~n448;
  assign po59 = ~n449 | ~n450;
  assign n452 = pi078 & po59;
  assign n453 = pi076 & n452;
  assign n454 = pi080 & n453;
  assign n455 = pi076 & pi077;
  assign n456 = pi078 & pi079;
  assign n457 = pi076 & n456;
  assign n458 = ~n454 & ~n455;
  assign n459 = ~pi097 & ~n457;
  assign po38 = ~n458 | ~n459;
  assign n461 = pi080 & n452;
  assign n462 = ~pi077 & ~n461;
  assign po39 = n456 | ~n462;
  assign n464 = pi080 & po59;
  assign po40 = pi079 | n464;
  assign n466 = pi120 & n443;
  assign n467 = ~pi117 & ~n466;
  assign po60 = n447 | ~n467;
  assign n469 = pi083 & po60;
  assign n470 = pi081 & n469;
  assign n471 = pi085 & n470;
  assign n472 = pi081 & pi082;
  assign n473 = pi083 & pi084;
  assign n474 = pi081 & n473;
  assign n475 = ~n471 & ~n472;
  assign n476 = ~pi098 & ~n474;
  assign po41 = ~n475 | ~n476;
  assign n478 = pi085 & n469;
  assign n479 = ~pi082 & ~n478;
  assign po42 = n473 | ~n479;
  assign n481 = pi085 & po60;
  assign po43 = pi084 | n481;
  assign n483 = pi095 & pi120;
  assign po61 = pi119 | n483;
  assign n485 = pi088 & po61;
  assign n486 = pi086 & n485;
  assign n487 = pi090 & n486;
  assign n488 = pi086 & pi087;
  assign n489 = pi088 & pi089;
  assign n490 = pi086 & n489;
  assign n491 = ~n487 & ~n488;
  assign n492 = ~pi099 & ~n490;
  assign po44 = ~n491 | ~n492;
  assign n494 = pi090 & n485;
  assign n495 = ~pi087 & ~n494;
  assign po45 = n489 | ~n495;
  assign n497 = pi090 & po61;
  assign po46 = pi089 | n497;
  assign n499 = pi093 & pi095;
  assign n500 = pi091 & n499;
  assign n501 = pi096 & n500;
  assign n502 = pi091 & pi092;
  assign n503 = pi093 & pi094;
  assign n504 = pi091 & n503;
  assign n505 = ~n501 & ~n502;
  assign n506 = ~pi100 & ~n504;
  assign po47 = ~n505 | ~n506;
  assign n508 = pi096 & n499;
  assign n509 = ~pi092 & ~n508;
  assign po48 = n503 | ~n509;
  assign n511 = pi095 & pi096;
  assign po49 = pi094 | n511;
endmodule



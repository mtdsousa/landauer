// Benchmark "i10" written by ABC on Sun Apr 22 21:43:04 2018

module i10 ( 
    pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008, pi009,
    pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018, pi019,
    pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028, pi029,
    pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038, pi039,
    pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048, pi049,
    pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058, pi059,
    pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068, pi069,
    pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078, pi079,
    pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088, pi089,
    pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098, pi099,
    pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109,
    pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118, pi119,
    pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128, pi129,
    pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138, pi139,
    pi140, pi141, pi142, pi143, pi144, pi145, pi146, pi147, pi148, pi149,
    pi150, pi151, pi152, pi153, pi154, pi155, pi156, pi157, pi158, pi159,
    pi160, pi161, pi162, pi163, pi164, pi165, pi166, pi167, pi168, pi169,
    pi170, pi171, pi172, pi173, pi174, pi175, pi176, pi177, pi178, pi179,
    pi180, pi181, pi182, pi183, pi184, pi185, pi186, pi187, pi188, pi189,
    pi190, pi191, pi192, pi193, pi194, pi195, pi196, pi197, pi198, pi199,
    pi200, pi201, pi202, pi203, pi204, pi205, pi206, pi207, pi208, pi209,
    pi210, pi211, pi212, pi213, pi214, pi215, pi216, pi217, pi218, pi219,
    pi220, pi221, pi222, pi223, pi224, pi225, pi226, pi227, pi228, pi229,
    pi230, pi231, pi232, pi233, pi234, pi235, pi236, pi237, pi238, pi239,
    pi240, pi241, pi242, pi243, pi244, pi245, pi246, pi247, pi248, pi249,
    pi250, pi251, pi252, pi253, pi254, pi255, pi256,
    po000, po001, po002, po003, po004, po005, po006, po007, po008, po009,
    po010, po011, po012, po013, po014, po015, po016, po017, po018, po019,
    po020, po021, po022, po023, po024, po025, po026, po027, po028, po029,
    po030, po031, po032, po033, po034, po035, po036, po037, po038, po039,
    po040, po041, po042, po043, po044, po045, po046, po047, po048, po049,
    po050, po051, po052, po053, po054, po055, po056, po057, po058, po059,
    po060, po061, po062, po063, po064, po065, po066, po067, po068, po069,
    po070, po071, po072, po073, po074, po075, po076, po077, po078, po079,
    po080, po081, po082, po083, po084, po085, po086, po087, po088, po089,
    po090, po091, po092, po093, po094, po095, po096, po097, po098, po099,
    po100, po101, po102, po103, po104, po105, po106, po107, po108, po109,
    po110, po111, po112, po113, po114, po115, po116, po117, po118, po119,
    po120, po121, po122, po123, po124, po125, po126, po127, po128, po129,
    po130, po131, po132, po133, po134, po135, po136, po137, po138, po139,
    po140, po141, po142, po143, po144, po145, po146, po147, po148, po149,
    po150, po151, po152, po153, po154, po155, po156, po157, po158, po159,
    po160, po161, po162, po163, po164, po165, po166, po167, po168, po169,
    po170, po171, po172, po173, po174, po175, po176, po177, po178, po179,
    po180, po181, po182, po183, po184, po185, po186, po187, po188, po189,
    po190, po191, po192, po193, po194, po195, po196, po197, po198, po199,
    po200, po201, po202, po203, po204, po205, po206, po207, po208, po209,
    po210, po211, po212, po213, po214, po215, po216, po217, po218, po219,
    po220, po221, po222, po223  );
  input  pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008,
    pi009, pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018,
    pi019, pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028,
    pi029, pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038,
    pi039, pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048,
    pi049, pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058,
    pi059, pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068,
    pi069, pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078,
    pi079, pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088,
    pi089, pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098,
    pi099, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108,
    pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118,
    pi119, pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128,
    pi129, pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138,
    pi139, pi140, pi141, pi142, pi143, pi144, pi145, pi146, pi147, pi148,
    pi149, pi150, pi151, pi152, pi153, pi154, pi155, pi156, pi157, pi158,
    pi159, pi160, pi161, pi162, pi163, pi164, pi165, pi166, pi167, pi168,
    pi169, pi170, pi171, pi172, pi173, pi174, pi175, pi176, pi177, pi178,
    pi179, pi180, pi181, pi182, pi183, pi184, pi185, pi186, pi187, pi188,
    pi189, pi190, pi191, pi192, pi193, pi194, pi195, pi196, pi197, pi198,
    pi199, pi200, pi201, pi202, pi203, pi204, pi205, pi206, pi207, pi208,
    pi209, pi210, pi211, pi212, pi213, pi214, pi215, pi216, pi217, pi218,
    pi219, pi220, pi221, pi222, pi223, pi224, pi225, pi226, pi227, pi228,
    pi229, pi230, pi231, pi232, pi233, pi234, pi235, pi236, pi237, pi238,
    pi239, pi240, pi241, pi242, pi243, pi244, pi245, pi246, pi247, pi248,
    pi249, pi250, pi251, pi252, pi253, pi254, pi255, pi256;
  output po000, po001, po002, po003, po004, po005, po006, po007, po008, po009,
    po010, po011, po012, po013, po014, po015, po016, po017, po018, po019,
    po020, po021, po022, po023, po024, po025, po026, po027, po028, po029,
    po030, po031, po032, po033, po034, po035, po036, po037, po038, po039,
    po040, po041, po042, po043, po044, po045, po046, po047, po048, po049,
    po050, po051, po052, po053, po054, po055, po056, po057, po058, po059,
    po060, po061, po062, po063, po064, po065, po066, po067, po068, po069,
    po070, po071, po072, po073, po074, po075, po076, po077, po078, po079,
    po080, po081, po082, po083, po084, po085, po086, po087, po088, po089,
    po090, po091, po092, po093, po094, po095, po096, po097, po098, po099,
    po100, po101, po102, po103, po104, po105, po106, po107, po108, po109,
    po110, po111, po112, po113, po114, po115, po116, po117, po118, po119,
    po120, po121, po122, po123, po124, po125, po126, po127, po128, po129,
    po130, po131, po132, po133, po134, po135, po136, po137, po138, po139,
    po140, po141, po142, po143, po144, po145, po146, po147, po148, po149,
    po150, po151, po152, po153, po154, po155, po156, po157, po158, po159,
    po160, po161, po162, po163, po164, po165, po166, po167, po168, po169,
    po170, po171, po172, po173, po174, po175, po176, po177, po178, po179,
    po180, po181, po182, po183, po184, po185, po186, po187, po188, po189,
    po190, po191, po192, po193, po194, po195, po196, po197, po198, po199,
    po200, po201, po202, po203, po204, po205, po206, po207, po208, po209,
    po210, po211, po212, po213, po214, po215, po216, po217, po218, po219,
    po220, po221, po222, po223;
  wire n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
    n493, n494, n495, n496, n497, n498, n499, n500, n502, n503, n504, n505,
    n506, n507, n508, n509, n510, n511, n512, n514, n515, n516, n517, n518,
    n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
    n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
    n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
    n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
    n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
    n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
    n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
    n603, n604, n605, n606, n608, n609, n610, n611, n612, n613, n614, n615,
    n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
    n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
    n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
    n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
    n664, n665, n666, n668, n669, n670, n671, n672, n673, n674, n675, n676,
    n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
    n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
    n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
    n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
    n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
    n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
    n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
    n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
    n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
    n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
    n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
    n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
    n822, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
    n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
    n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
    n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
    n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
    n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
    n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n908,
    n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
    n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
    n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
    n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
    n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
    n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
    n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
    n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
    n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
    n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
    n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
    n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
    n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
    n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
    n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
    n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
    n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
    n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
    n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
    n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
    n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
    n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
    n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
    n1154, n1155, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
    n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
    n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
    n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
    n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
    n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
    n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
    n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
    n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
    n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
    n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
    n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
    n1275, n1276, n1279, n1280, n1281, n1289, n1293, n1294, n1295, n1296,
    n1297, n1298, n1299, n1300, n1302, n1303, n1304, n1305, n1307, n1308,
    n1309, n1310, n1311, n1312, n1314, n1315, n1316, n1317, n1318, n1319,
    n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
    n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
    n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
    n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359,
    n1360, n1361, n1362, n1364, n1365, n1366, n1367, n1368, n1369, n1370,
    n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380,
    n1381, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391,
    n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1402,
    n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
    n1413, n1414, n1415, n1416, n1417, n1419, n1420, n1421, n1422, n1423,
    n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433,
    n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443,
    n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453,
    n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464,
    n1465, n1466, n1467, n1468, n1470, n1471, n1472, n1473, n1474, n1475,
    n1477, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487,
    n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497,
    n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507,
    n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517,
    n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527,
    n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537,
    n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547,
    n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557,
    n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567,
    n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577,
    n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587,
    n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597,
    n1598, n1599, n1600, n1602, n1603, n1604, n1605, n1606, n1607, n1608,
    n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1619, n1620, n1621,
    n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631,
    n1633, n1635, n1636, n1637, n1638, n1639, n1640, n1642, n1643, n1644,
    n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654,
    n1655, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669,
    n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1681,
    n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691,
    n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701,
    n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713,
    n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723,
    n1724, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735,
    n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745,
    n1746, n1747, n1748, n1749, n1750, n1753, n1754, n1755, n1756, n1757,
    n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767,
    n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1779,
    n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789,
    n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799,
    n1800, n1801, n1802, n1805, n1806, n1807, n1808, n1809, n1810, n1811,
    n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821,
    n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1832, n1833,
    n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843,
    n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853,
    n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865,
    n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1876,
    n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1887,
    n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897,
    n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908,
    n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918,
    n1919, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929,
    n1930, n1931, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940,
    n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950,
    n1951, n1952, n1953, n1955, n1956, n1957, n1958, n1959, n1960, n1961,
    n1962, n1963, n1964, n1965, n1966, n1968, n1969, n1970, n1971, n1972,
    n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
    n1983, n1984, n1985, n1986, n1987, n1988, n1990, n1991, n1992, n1993,
    n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2003, n2004,
    n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014,
    n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024,
    n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034,
    n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2044, n2045,
    n2046, n2047, n2048, n2050, n2051, n2052, n2053, n2054, n2055, n2056,
    n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066,
    n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076,
    n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086,
    n2087, n2088, n2089, n2091, n2092, n2093, n2094, n2095, n2097, n2098,
    n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108,
    n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118,
    n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128,
    n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2139,
    n2140, n2141, n2142, n2143, n2145, n2146, n2147, n2148, n2149, n2150,
    n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2161,
    n2163, n2164, n2165, n2166, n2168, n2169, n2170, n2171, n2173, n2174,
    n2175, n2176, n2178, n2179, n2180, n2181, n2183, n2184, n2185, n2186,
    n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2195, n2196, n2197,
    n2199, n2200, n2202, n2203, n2204, n2206, n2207, n2208, n2209, n2210,
    n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220,
    n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230,
    n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240,
    n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250,
    n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2259, n2261, n2262,
    n2263, n2264, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276,
    n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286,
    n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296,
    n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306,
    n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316,
    n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326,
    n2327, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337,
    n2338, n2339, n2342, n2343, n2344, n2346, n2347, n2348, n2349, n2350,
    n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361,
    n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
    n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384,
    n2385, n2386, n2387, n2388, n2397, n2398, n2399, n2400, n2401, n2402,
    n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
    n2413, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423,
    n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433,
    n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2443, n2444,
    n2445, n2446, n2447, n2449, n2450, n2451, n2452, n2453, n2455, n2456,
    n2457, n2458, n2459, n2461, n2462, n2463, n2464, n2465, n2467, n2468,
    n2469, n2470, n2471, n2473, n2474, n2475, n2476, n2477, n2478, n2479,
    n2481, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491,
    n2492, n2493, n2494, n2495, n2496, n2498, n2499, n2500, n2502, n2503,
    n2504, n2505, n2507, n2508, n2509, n2510, n2512, n2513, n2514, n2515,
    n2516, n2517, n2518, n2519, n2520, n2525, n2527, n2528, n2531, n2532,
    n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2542, n2543,
    n2544, n2545, n2546, n2547, n2548, n2550, n2551, n2552, n2553, n2554,
    n2555, n2556, n2558, n2559, n2561, n2562, n2563, n2564, n2566, n2567,
    n2568, n2569, n2570, n2571, n2572, n2574, n2575, n2576, n2577, n2578,
    n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588,
    n2589, n2590, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599,
    n2600, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610,
    n2611, n2612, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621,
    n2622, n2624, n2626, n2627, n2629, n2630, n2631, n2632, n2633, n2634,
    n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2645, n2646,
    n2648, n2649, n2650, n2651, n2652, n2653, n2655, n2656, n2657, n2658,
    n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668,
    n2669, n2670, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679,
    n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689,
    n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700,
    n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710,
    n2711, n2712, n2713, n2714, n2716, n2717, n2718, n2719, n2720, n2721,
    n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731,
    n2732, n2733, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
    n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
    n2753, n2754, n2755, n2757, n2758, n2759, n2760, n2761, n2762, n2763,
    n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773,
    n2774, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2785,
    n2786, n2787, n2788, n2790, n2791, n2792, n2793, n2795, n2796, n2797,
    n2798, n2799, n2800, n2801, n2802, n2803, n2805, n2806, n2807, n2808,
    n2809, n2810, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819,
    n2820, n2821, n2822, n2823, n2825, n2826, n2827, n2828, n2829, n2830,
    n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2842,
    n2843, n2844, n2845, n2846, n2847, n2849, n2850, n2851, n2852, n2853,
    n2854, n2855, n2856, n2858, n2859, n2860, n2861, n2862, n2864, n2865,
    n2866, n2867, n2868, n2869, n2870, n2872, n2873, n2875, n2876, n2877,
    n2878, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888,
    n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898,
    n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2908, n2909, n2910,
    n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920,
    n2921, n2922, n2924, n2925, n2926, n2927, n2928, n2930, n2931, n2932,
    n2933, n2934, n2936, n2937, n2938, n2939, n2940, n2942, n2943, n2944,
    n2945, n2946, n2948, n2949, n2950, n2951, n2952, n2954, n2955, n2956,
    n2957, n2958, n2959, n2960, n2961, n2963, n2964, n2965, n2966, n2968,
    n2969, n2971, n2972, n2974, n2976, n2977, n2978, n2979, n2980, n2981,
    n2983, n2984, n2985, n2986, n2988, n2989, n2990, n2991, n2993, n2994,
    n2995, n2996, n2998, n2999, n3000, n3001, n3003, n3004, n3005, n3006,
    n3008, n3009, n3010, n3011, n3013, n3014, n3015, n3016, n3018, n3019,
    n3020, n3021, n3023, n3024, n3025, n3026, n3028, n3029, n3030, n3031,
    n3033, n3034, n3035, n3036, n3038, n3039, n3040, n3041, n3043, n3044,
    n3045, n3046, n3048, n3049, n3051, n3052, n3053, n3054, n3056, n3057,
    n3058, n3060, n3061, n3063, n3064, n3066, n3067, n3069, n3071, n3073,
    n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3083, n3084,
    n3085, n3086, n3087, n3088, n3089, n3090, n3092, n3093, n3094, n3095,
    n3096, n3097, n3098, n3099, n3100, n3102, n3103, n3104, n3105, n3106,
    n3107, n3108, n3109, n3111, n3112, n3113, n3114, n3115, n3117, n3118,
    n3119, n3120, n3122, n3123, n3124, n3125, n3127, n3128, n3129, n3131,
    n3132, n3133, n3135, n3136, n3138, n3139, n3141, n3142, n3143, n3144,
    n3146, n3147, n3148, n3150, n3151, n3152, n3154, n3155;
  assign n482 = pi029 & ~pi053;
  assign n483 = pi054 & n482;
  assign n484 = pi055 & n483;
  assign n485 = ~pi056 & n484;
  assign n486 = ~pi053 & ~pi055;
  assign n487 = ~pi054 & n486;
  assign n488 = pi054 & ~pi055;
  assign n489 = ~pi053 & n488;
  assign n490 = pi026 & pi028;
  assign n491 = ~pi056 & n490;
  assign n492 = n489 & n491;
  assign n493 = pi029 & n492;
  assign n494 = pi027 & n493;
  assign n495 = ~pi026 & pi028;
  assign n496 = ~pi056 & n495;
  assign n497 = n489 & n496;
  assign n498 = pi029 & n497;
  assign n499 = pi027 & n498;
  assign n500 = ~n494 & ~n499;
  assign po065 = pi069 | pi076;
  assign n502 = ~pi067 & ~n500;
  assign n503 = ~po065 & n502;
  assign n504 = ~n485 & ~n487;
  assign n505 = ~n503 & n504;
  assign n506 = pi019 & ~pi061;
  assign n507 = pi075 & n506;
  assign n508 = ~pi060 & n507;
  assign n509 = ~pi062 & n508;
  assign n510 = pi068 & ~n505;
  assign n511 = ~pi183 & n510;
  assign n512 = ~n509 & n511;
  assign po052 = ~pi182 & n512;
  assign n514 = pi019 & pi063;
  assign n515 = pi191 & n514;
  assign n516 = pi061 & n515;
  assign n517 = pi075 & n516;
  assign n518 = pi060 & n517;
  assign n519 = pi062 & n518;
  assign n520 = pi058 & n519;
  assign n521 = pi064 & n520;
  assign n522 = pi059 & n521;
  assign n523 = po052 & n522;
  assign n524 = pi062 & pi063;
  assign n525 = pi061 & n524;
  assign n526 = pi075 & n525;
  assign n527 = pi060 & n526;
  assign n528 = pi191 & n527;
  assign n529 = ~pi189 & n528;
  assign n530 = pi058 & n529;
  assign n531 = pi064 & n530;
  assign n532 = pi059 & n531;
  assign n533 = ~n523 & ~n532;
  assign n534 = ~pi192 & n533;
  assign n535 = pi055 & pi056;
  assign n536 = pi054 & n535;
  assign n537 = ~pi053 & n536;
  assign n538 = ~pi016 & n485;
  assign n539 = pi167 & n538;
  assign n540 = pi168 & ~n539;
  assign n541 = n537 & ~n540;
  assign n542 = ~pi015 & n541;
  assign n543 = ~pi054 & pi055;
  assign n544 = ~pi053 & n543;
  assign n545 = ~n487 & ~n544;
  assign n546 = ~pi029 & ~pi053;
  assign n547 = pi054 & n546;
  assign n548 = pi055 & n547;
  assign n549 = ~pi056 & n548;
  assign n550 = ~n538 & n545;
  assign n551 = ~n549 & n550;
  assign n552 = ~pi016 & ~n551;
  assign n553 = n537 & n540;
  assign n554 = ~pi015 & ~pi163;
  assign n555 = n541 & ~n554;
  assign n556 = ~n552 & ~n553;
  assign n557 = ~n555 & n556;
  assign n558 = pi045 & ~n534;
  assign n559 = ~n542 & n558;
  assign n560 = n557 & n559;
  assign n561 = ~pi015 & pi029;
  assign n562 = ~n540 & n561;
  assign n563 = n537 & n562;
  assign n564 = n534 & n563;
  assign n565 = n557 & n564;
  assign n566 = ~n537 & ~n538;
  assign n567 = ~n549 & n566;
  assign n568 = pi118 & ~n545;
  assign n569 = n567 & n568;
  assign n570 = pi128 & n545;
  assign n571 = ~n567 & n570;
  assign n572 = ~n569 & ~n571;
  assign n573 = n534 & ~n572;
  assign n574 = ~n542 & n573;
  assign n575 = ~n557 & n574;
  assign n576 = ~n560 & ~n565;
  assign n577 = ~n575 & n576;
  assign n578 = po052 & n534;
  assign n579 = ~n577 & ~n578;
  assign n580 = ~n578 & n579;
  assign n581 = ~pi004 & ~pi015;
  assign n582 = ~pi163 & n581;
  assign n583 = po052 & ~n582;
  assign n584 = pi002 & n583;
  assign n585 = pi133 & ~n583;
  assign n586 = ~n583 & n585;
  assign n587 = ~n584 & ~n586;
  assign n588 = n578 & ~n587;
  assign n589 = n578 & n588;
  assign n590 = ~n580 & ~n589;
  assign n591 = pi056 & n544;
  assign n592 = ~n538 & ~n591;
  assign n593 = pi163 & ~n592;
  assign n594 = pi026 & ~pi028;
  assign n595 = ~pi056 & n594;
  assign n596 = n489 & n595;
  assign n597 = pi029 & n596;
  assign n598 = pi027 & n597;
  assign n599 = ~pi016 & n487;
  assign n600 = ~pi029 & ~pi056;
  assign n601 = n599 & n600;
  assign n602 = pi028 & n601;
  assign n603 = pi065 & n602;
  assign n604 = ~pi066 & n603;
  assign n605 = ~pi065 & n602;
  assign n606 = ~pi066 & n605;
  assign po051 = ~pi056 & n599;
  assign n608 = ~pi028 & ~pi029;
  assign n609 = po051 & n608;
  assign n610 = pi065 & n609;
  assign n611 = ~pi066 & n610;
  assign n612 = pi028 & po051;
  assign n613 = pi029 & n612;
  assign n614 = ~pi028 & po051;
  assign n615 = pi029 & n614;
  assign n616 = ~pi065 & n609;
  assign n617 = pi066 & n616;
  assign n618 = pi066 & n610;
  assign n619 = pi066 & n605;
  assign n620 = ~n611 & ~n613;
  assign n621 = ~n604 & ~n606;
  assign n622 = n620 & n621;
  assign n623 = ~n618 & ~n619;
  assign n624 = ~n615 & ~n617;
  assign n625 = n623 & n624;
  assign n626 = n622 & n625;
  assign n627 = pi057 & ~n545;
  assign n628 = ~n626 & n627;
  assign n629 = pi163 & n628;
  assign n630 = pi056 & n599;
  assign n631 = n627 & n630;
  assign n632 = pi163 & n631;
  assign n633 = pi004 & n631;
  assign n634 = pi004 & n628;
  assign n635 = ~n633 & ~n634;
  assign n636 = ~n629 & ~n632;
  assign n637 = n635 & n636;
  assign n638 = n538 & ~n540;
  assign n639 = ~pi028 & ~pi056;
  assign n640 = n544 & n639;
  assign n641 = pi029 & n640;
  assign n642 = ~pi029 & n640;
  assign n643 = pi028 & ~pi056;
  assign n644 = n544 & n643;
  assign n645 = ~pi029 & n644;
  assign n646 = ~n641 & ~n642;
  assign n647 = ~n645 & n646;
  assign n648 = ~n591 & n626;
  assign n649 = ~n638 & n647;
  assign n650 = ~n630 & n649;
  assign n651 = n648 & n650;
  assign n652 = ~pi004 & ~pi164;
  assign n653 = ~pi165 & n652;
  assign n654 = n637 & ~n651;
  assign n655 = ~n653 & n654;
  assign n656 = n534 & ~n549;
  assign n657 = ~n537 & n656;
  assign n658 = pi164 & n657;
  assign n659 = ~pi004 & n658;
  assign n660 = ~n598 & ~n655;
  assign n661 = ~n659 & n660;
  assign n662 = ~n593 & ~n661;
  assign n663 = ~n590 & ~n662;
  assign n664 = n661 & n663;
  assign n665 = pi147 & n662;
  assign n666 = ~n661 & n665;
  assign po000 = ~n664 & ~n666;
  assign n668 = ~pi026 & ~pi028;
  assign n669 = pi056 & n668;
  assign n670 = n489 & n669;
  assign n671 = ~pi029 & n670;
  assign n672 = ~pi027 & n671;
  assign n673 = ~po065 & n672;
  assign n674 = n534 & ~n673;
  assign n675 = ~pi083 & pi207;
  assign n676 = ~pi082 & pi208;
  assign n677 = ~pi081 & pi209;
  assign n678 = ~pi010 & pi011;
  assign n679 = n677 & n678;
  assign n680 = ~n677 & ~n678;
  assign n681 = ~n679 & ~n680;
  assign n682 = n676 & n681;
  assign n683 = ~n676 & ~n681;
  assign n684 = ~n682 & ~n683;
  assign n685 = n675 & n684;
  assign n686 = ~n675 & ~n684;
  assign n687 = ~n685 & ~n686;
  assign n688 = n675 & ~n687;
  assign n689 = n675 & n688;
  assign n690 = pi083 & ~pi207;
  assign n691 = ~n687 & n690;
  assign n692 = n690 & n691;
  assign n693 = ~n687 & ~n690;
  assign n694 = ~n690 & n693;
  assign n695 = ~n692 & ~n694;
  assign n696 = ~n675 & n695;
  assign n697 = ~n675 & n696;
  assign n698 = ~n689 & ~n697;
  assign n699 = pi093 & ~n545;
  assign n700 = n567 & n699;
  assign n701 = pi105 & n545;
  assign n702 = ~n567 & n701;
  assign n703 = ~n700 & ~n702;
  assign n704 = ~n557 & ~n578;
  assign n705 = ~n703 & n704;
  assign n706 = n534 & n705;
  assign n707 = ~n542 & n706;
  assign n708 = ~n578 & n707;
  assign n709 = ~n662 & n708;
  assign n710 = n661 & n709;
  assign n711 = pi003 & n662;
  assign n712 = ~n661 & n711;
  assign po078 = n710 | n712;
  assign n714 = ~n698 & ~po078;
  assign n715 = n698 & po078;
  assign n716 = ~n714 & ~n715;
  assign n717 = pi082 & ~pi208;
  assign n718 = pi081 & ~pi209;
  assign n719 = pi010 & ~pi011;
  assign n720 = ~n678 & ~n719;
  assign n721 = n718 & ~n720;
  assign n722 = ~n718 & n720;
  assign n723 = ~n721 & ~n722;
  assign n724 = n677 & ~n678;
  assign n725 = ~n723 & ~n724;
  assign n726 = n723 & n724;
  assign n727 = ~n725 & ~n726;
  assign n728 = n717 & n727;
  assign n729 = ~n717 & ~n727;
  assign n730 = ~n728 & ~n729;
  assign n731 = n676 & ~n681;
  assign n732 = ~n730 & ~n731;
  assign n733 = n730 & n731;
  assign n734 = ~n732 & ~n733;
  assign n735 = n690 & ~n734;
  assign n736 = n675 & ~n684;
  assign n737 = n690 & n736;
  assign n738 = ~n734 & n736;
  assign n739 = ~n735 & ~n737;
  assign n740 = ~n738 & n739;
  assign n741 = pi083 & pi207;
  assign n742 = n717 & ~n727;
  assign n743 = n717 & n731;
  assign n744 = ~n727 & n731;
  assign n745 = ~n742 & ~n743;
  assign n746 = ~n744 & n745;
  assign n747 = pi082 & pi208;
  assign n748 = n718 & n720;
  assign n749 = n718 & n724;
  assign n750 = n720 & n724;
  assign n751 = ~n748 & ~n749;
  assign n752 = ~n750 & n751;
  assign n753 = pi081 & pi209;
  assign n754 = ~pi010 & ~pi011;
  assign n755 = n753 & ~n754;
  assign n756 = ~n753 & n754;
  assign n757 = ~n755 & ~n756;
  assign n758 = ~n752 & n757;
  assign n759 = n752 & ~n757;
  assign n760 = ~n758 & ~n759;
  assign n761 = n747 & n760;
  assign n762 = ~n747 & ~n760;
  assign n763 = ~n761 & ~n762;
  assign n764 = ~n746 & n763;
  assign n765 = n746 & ~n763;
  assign n766 = ~n764 & ~n765;
  assign n767 = n741 & n766;
  assign n768 = ~n741 & ~n766;
  assign n769 = ~n767 & ~n768;
  assign n770 = ~n740 & n769;
  assign n771 = n740 & ~n769;
  assign n772 = ~n770 & ~n771;
  assign n773 = n675 & ~n772;
  assign n774 = n675 & n773;
  assign n775 = n690 & ~n772;
  assign n776 = n690 & n775;
  assign n777 = n690 & n734;
  assign n778 = ~n690 & ~n734;
  assign n779 = ~n777 & ~n778;
  assign n780 = ~n736 & ~n779;
  assign n781 = n736 & n779;
  assign n782 = ~n780 & ~n781;
  assign n783 = n687 & n782;
  assign n784 = ~n772 & ~n783;
  assign n785 = n772 & n783;
  assign n786 = ~n784 & ~n785;
  assign n787 = ~n687 & ~n782;
  assign n788 = ~n783 & ~n787;
  assign n789 = ~n687 & n788;
  assign n790 = ~n786 & ~n789;
  assign n791 = n786 & n789;
  assign n792 = ~n790 & ~n791;
  assign n793 = ~n690 & ~n792;
  assign n794 = ~n690 & n793;
  assign n795 = ~n776 & ~n794;
  assign n796 = n690 & ~n782;
  assign n797 = n690 & n796;
  assign n798 = n687 & ~n788;
  assign n799 = ~n789 & ~n798;
  assign n800 = ~n690 & ~n799;
  assign n801 = ~n690 & n800;
  assign n802 = ~n797 & ~n801;
  assign n803 = n695 & n802;
  assign n804 = ~n795 & ~n803;
  assign n805 = n795 & n803;
  assign n806 = ~n804 & ~n805;
  assign n807 = ~n675 & ~n806;
  assign n808 = ~n675 & n807;
  assign n809 = ~n774 & ~n808;
  assign n810 = pi095 & ~n545;
  assign n811 = n567 & n810;
  assign n812 = pi107 & n545;
  assign n813 = ~n567 & n812;
  assign n814 = ~n811 & ~n813;
  assign n815 = n704 & ~n814;
  assign n816 = n534 & n815;
  assign n817 = ~n542 & n816;
  assign n818 = ~n578 & n817;
  assign n819 = ~n662 & n818;
  assign n820 = n661 & n819;
  assign n821 = pi001 & n662;
  assign n822 = ~n661 & n821;
  assign po080 = n820 | n822;
  assign n824 = ~n809 & ~po080;
  assign n825 = n809 & po080;
  assign n826 = ~n824 & ~n825;
  assign n827 = n753 & n754;
  assign n828 = ~n752 & n753;
  assign n829 = ~n752 & n754;
  assign n830 = ~n827 & ~n828;
  assign n831 = ~n829 & n830;
  assign n832 = n754 & n831;
  assign n833 = ~n754 & ~n831;
  assign n834 = ~n832 & ~n833;
  assign n835 = n747 & ~n760;
  assign n836 = ~n746 & n747;
  assign n837 = ~n746 & ~n760;
  assign n838 = ~n835 & ~n836;
  assign n839 = ~n837 & n838;
  assign n840 = ~n834 & n839;
  assign n841 = n834 & ~n839;
  assign n842 = ~n840 & ~n841;
  assign n843 = n741 & ~n766;
  assign n844 = ~n740 & n741;
  assign n845 = ~n740 & ~n766;
  assign n846 = ~n843 & ~n844;
  assign n847 = ~n845 & n846;
  assign n848 = ~n842 & n847;
  assign n849 = n842 & ~n847;
  assign n850 = ~n848 & ~n849;
  assign n851 = n675 & ~n850;
  assign n852 = n675 & n851;
  assign n853 = n690 & ~n850;
  assign n854 = n690 & n853;
  assign n855 = ~n785 & ~n850;
  assign n856 = n785 & n850;
  assign n857 = ~n855 & ~n856;
  assign n858 = ~n791 & ~n857;
  assign n859 = n791 & n857;
  assign n860 = ~n858 & ~n859;
  assign n861 = ~n690 & ~n860;
  assign n862 = ~n690 & n861;
  assign n863 = ~n854 & ~n862;
  assign n864 = ~n805 & ~n863;
  assign n865 = n805 & n863;
  assign n866 = ~n864 & ~n865;
  assign n867 = ~n675 & ~n866;
  assign n868 = ~n675 & n867;
  assign n869 = ~n852 & ~n868;
  assign n870 = pi096 & ~n545;
  assign n871 = n567 & n870;
  assign n872 = pi108 & n545;
  assign n873 = ~n567 & n872;
  assign n874 = ~n871 & ~n873;
  assign n875 = n704 & ~n874;
  assign n876 = n534 & n875;
  assign n877 = ~n542 & n876;
  assign n878 = ~n578 & n877;
  assign n879 = ~n662 & n878;
  assign n880 = n661 & n879;
  assign n881 = pi000 & n662;
  assign n882 = ~n661 & n881;
  assign po081 = n880 | n882;
  assign n884 = ~n869 & ~po081;
  assign n885 = n869 & po081;
  assign n886 = ~n884 & ~n885;
  assign n887 = n675 & ~n782;
  assign n888 = n675 & n887;
  assign n889 = ~n695 & ~n802;
  assign n890 = ~n803 & ~n889;
  assign n891 = ~n675 & ~n890;
  assign n892 = ~n675 & n891;
  assign n893 = ~n888 & ~n892;
  assign n894 = pi094 & ~n545;
  assign n895 = n567 & n894;
  assign n896 = pi106 & n545;
  assign n897 = ~n567 & n896;
  assign n898 = ~n895 & ~n897;
  assign n899 = n704 & ~n898;
  assign n900 = n534 & n899;
  assign n901 = ~n542 & n900;
  assign n902 = ~n578 & n901;
  assign n903 = ~n662 & n902;
  assign n904 = n661 & n903;
  assign n905 = pi002 & n662;
  assign n906 = ~n661 & n905;
  assign po079 = n904 | n906;
  assign n908 = ~n893 & ~po079;
  assign n909 = n893 & po079;
  assign n910 = ~n908 & ~n909;
  assign n911 = ~pi083 & ~pi207;
  assign n912 = ~n673 & n716;
  assign n913 = n826 & n912;
  assign n914 = n886 & n913;
  assign n915 = n910 & n914;
  assign n916 = ~n911 & n915;
  assign n917 = n676 & ~n684;
  assign n918 = n676 & n917;
  assign n919 = ~n684 & n717;
  assign n920 = n717 & n919;
  assign n921 = ~n684 & ~n717;
  assign n922 = ~n717 & n921;
  assign n923 = ~n920 & ~n922;
  assign n924 = ~n676 & n923;
  assign n925 = ~n676 & n924;
  assign n926 = ~n918 & ~n925;
  assign n927 = ~po078 & ~n926;
  assign n928 = po078 & n926;
  assign n929 = ~n927 & ~n928;
  assign n930 = n676 & ~n766;
  assign n931 = n676 & n930;
  assign n932 = n717 & ~n766;
  assign n933 = n717 & n932;
  assign n934 = n684 & n734;
  assign n935 = ~n766 & ~n934;
  assign n936 = n766 & n934;
  assign n937 = ~n935 & ~n936;
  assign n938 = ~n684 & ~n734;
  assign n939 = ~n934 & ~n938;
  assign n940 = ~n684 & n939;
  assign n941 = ~n937 & ~n940;
  assign n942 = n937 & n940;
  assign n943 = ~n941 & ~n942;
  assign n944 = ~n717 & ~n943;
  assign n945 = ~n717 & n944;
  assign n946 = ~n933 & ~n945;
  assign n947 = n717 & ~n734;
  assign n948 = n717 & n947;
  assign n949 = n684 & ~n939;
  assign n950 = ~n940 & ~n949;
  assign n951 = ~n717 & ~n950;
  assign n952 = ~n717 & n951;
  assign n953 = ~n948 & ~n952;
  assign n954 = n923 & n953;
  assign n955 = ~n946 & ~n954;
  assign n956 = n946 & n954;
  assign n957 = ~n955 & ~n956;
  assign n958 = ~n676 & ~n957;
  assign n959 = ~n676 & n958;
  assign n960 = ~n931 & ~n959;
  assign n961 = ~po080 & ~n960;
  assign n962 = po080 & n960;
  assign n963 = ~n961 & ~n962;
  assign n964 = n676 & ~n842;
  assign n965 = n676 & n964;
  assign n966 = n717 & ~n842;
  assign n967 = n717 & n966;
  assign n968 = ~n842 & ~n936;
  assign n969 = n842 & n936;
  assign n970 = ~n968 & ~n969;
  assign n971 = ~n942 & ~n970;
  assign n972 = n942 & n970;
  assign n973 = ~n971 & ~n972;
  assign n974 = ~n717 & ~n973;
  assign n975 = ~n717 & n974;
  assign n976 = ~n967 & ~n975;
  assign n977 = ~n956 & ~n976;
  assign n978 = n956 & n976;
  assign n979 = ~n977 & ~n978;
  assign n980 = ~n676 & ~n979;
  assign n981 = ~n676 & n980;
  assign n982 = ~n965 & ~n981;
  assign n983 = ~po081 & ~n982;
  assign n984 = po081 & n982;
  assign n985 = ~n983 & ~n984;
  assign n986 = n676 & ~n734;
  assign n987 = n676 & n986;
  assign n988 = ~n923 & ~n953;
  assign n989 = ~n954 & ~n988;
  assign n990 = ~n676 & ~n989;
  assign n991 = ~n676 & n990;
  assign n992 = ~n987 & ~n991;
  assign n993 = ~po079 & ~n992;
  assign n994 = po079 & n992;
  assign n995 = ~n993 & ~n994;
  assign n996 = ~pi082 & ~pi208;
  assign n997 = ~n673 & n929;
  assign n998 = n963 & n997;
  assign n999 = n985 & n998;
  assign n1000 = n995 & n999;
  assign n1001 = ~n996 & n1000;
  assign n1002 = n677 & ~n681;
  assign n1003 = n677 & n1002;
  assign n1004 = ~n681 & n718;
  assign n1005 = n718 & n1004;
  assign n1006 = ~n681 & ~n718;
  assign n1007 = ~n718 & n1006;
  assign n1008 = ~n1005 & ~n1007;
  assign n1009 = ~n677 & n1008;
  assign n1010 = ~n677 & n1009;
  assign n1011 = ~n1003 & ~n1010;
  assign n1012 = ~po078 & ~n1011;
  assign n1013 = po078 & n1011;
  assign n1014 = ~n1012 & ~n1013;
  assign n1015 = n677 & ~n760;
  assign n1016 = n677 & n1015;
  assign n1017 = n718 & ~n760;
  assign n1018 = n718 & n1017;
  assign n1019 = n681 & n727;
  assign n1020 = ~n760 & ~n1019;
  assign n1021 = n760 & n1019;
  assign n1022 = ~n1020 & ~n1021;
  assign n1023 = ~n681 & ~n727;
  assign n1024 = ~n1019 & ~n1023;
  assign n1025 = ~n681 & n1024;
  assign n1026 = ~n1022 & ~n1025;
  assign n1027 = n1022 & n1025;
  assign n1028 = ~n1026 & ~n1027;
  assign n1029 = ~n718 & ~n1028;
  assign n1030 = ~n718 & n1029;
  assign n1031 = ~n1018 & ~n1030;
  assign n1032 = n718 & ~n727;
  assign n1033 = n718 & n1032;
  assign n1034 = n681 & ~n1024;
  assign n1035 = ~n1025 & ~n1034;
  assign n1036 = ~n718 & ~n1035;
  assign n1037 = ~n718 & n1036;
  assign n1038 = ~n1033 & ~n1037;
  assign n1039 = n1008 & n1038;
  assign n1040 = ~n1031 & ~n1039;
  assign n1041 = n1031 & n1039;
  assign n1042 = ~n1040 & ~n1041;
  assign n1043 = ~n677 & ~n1042;
  assign n1044 = ~n677 & n1043;
  assign n1045 = ~n1016 & ~n1044;
  assign n1046 = ~po080 & ~n1045;
  assign n1047 = po080 & n1045;
  assign n1048 = ~n1046 & ~n1047;
  assign n1049 = n677 & ~n834;
  assign n1050 = n677 & n1049;
  assign n1051 = n718 & ~n834;
  assign n1052 = n718 & n1051;
  assign n1053 = ~n834 & ~n1021;
  assign n1054 = n834 & n1021;
  assign n1055 = ~n1053 & ~n1054;
  assign n1056 = ~n1027 & ~n1055;
  assign n1057 = n1027 & n1055;
  assign n1058 = ~n1056 & ~n1057;
  assign n1059 = ~n718 & ~n1058;
  assign n1060 = ~n718 & n1059;
  assign n1061 = ~n1052 & ~n1060;
  assign n1062 = ~n1041 & ~n1061;
  assign n1063 = n1041 & n1061;
  assign n1064 = ~n1062 & ~n1063;
  assign n1065 = ~n677 & ~n1064;
  assign n1066 = ~n677 & n1065;
  assign n1067 = ~n1050 & ~n1066;
  assign n1068 = ~po081 & ~n1067;
  assign n1069 = po081 & n1067;
  assign n1070 = ~n1068 & ~n1069;
  assign n1071 = n677 & ~n727;
  assign n1072 = n677 & n1071;
  assign n1073 = ~n1008 & ~n1038;
  assign n1074 = ~n1039 & ~n1073;
  assign n1075 = ~n677 & ~n1074;
  assign n1076 = ~n677 & n1075;
  assign n1077 = ~n1072 & ~n1076;
  assign n1078 = ~po079 & ~n1077;
  assign n1079 = po079 & n1077;
  assign n1080 = ~n1078 & ~n1079;
  assign n1081 = ~pi081 & ~pi209;
  assign n1082 = ~n673 & n1014;
  assign n1083 = n1048 & n1082;
  assign n1084 = n1070 & n1083;
  assign n1085 = n1080 & n1084;
  assign n1086 = ~n1081 & n1085;
  assign n1087 = ~n673 & ~po078;
  assign n1088 = ~po080 & n1087;
  assign n1089 = ~po081 & n1088;
  assign n1090 = ~po079 & n1089;
  assign n1091 = ~n754 & n1090;
  assign n1092 = ~n673 & po079;
  assign n1093 = ~po080 & n1092;
  assign n1094 = ~po081 & n1093;
  assign n1095 = ~po078 & n1094;
  assign n1096 = pi010 & n1095;
  assign n1097 = pi011 & n1096;
  assign n1098 = n681 & ~po078;
  assign n1099 = ~n681 & po078;
  assign n1100 = ~n1098 & ~n1099;
  assign n1101 = ~po080 & ~n1022;
  assign n1102 = po080 & n1022;
  assign n1103 = ~n1101 & ~n1102;
  assign n1104 = ~po081 & ~n1055;
  assign n1105 = po081 & n1055;
  assign n1106 = ~n1104 & ~n1105;
  assign n1107 = ~po079 & ~n1024;
  assign n1108 = po079 & n1024;
  assign n1109 = ~n1107 & ~n1108;
  assign n1110 = ~n673 & n1100;
  assign n1111 = n1103 & n1110;
  assign n1112 = n1106 & n1111;
  assign n1113 = n1109 & n1112;
  assign n1114 = n753 & n1113;
  assign n1115 = n684 & ~po078;
  assign n1116 = ~n684 & po078;
  assign n1117 = ~n1115 & ~n1116;
  assign n1118 = ~po080 & ~n937;
  assign n1119 = po080 & n937;
  assign n1120 = ~n1118 & ~n1119;
  assign n1121 = ~po081 & ~n970;
  assign n1122 = po081 & n970;
  assign n1123 = ~n1121 & ~n1122;
  assign n1124 = ~po079 & ~n939;
  assign n1125 = po079 & n939;
  assign n1126 = ~n1124 & ~n1125;
  assign n1127 = ~n673 & n1117;
  assign n1128 = n1120 & n1127;
  assign n1129 = n1123 & n1128;
  assign n1130 = n1126 & n1129;
  assign n1131 = n747 & n1130;
  assign n1132 = n687 & ~po078;
  assign n1133 = ~n687 & po078;
  assign n1134 = ~n1132 & ~n1133;
  assign n1135 = ~n786 & ~po080;
  assign n1136 = n786 & po080;
  assign n1137 = ~n1135 & ~n1136;
  assign n1138 = ~n857 & ~po081;
  assign n1139 = n857 & po081;
  assign n1140 = ~n1138 & ~n1139;
  assign n1141 = ~n788 & ~po079;
  assign n1142 = n788 & po079;
  assign n1143 = ~n1141 & ~n1142;
  assign n1144 = ~n673 & n1134;
  assign n1145 = n1137 & n1144;
  assign n1146 = n1140 & n1145;
  assign n1147 = n1143 & n1146;
  assign n1148 = n741 & n1147;
  assign n1149 = n674 & ~n916;
  assign n1150 = ~n1001 & n1149;
  assign n1151 = ~n1086 & n1150;
  assign n1152 = ~n1091 & n1151;
  assign n1153 = ~n1097 & n1152;
  assign n1154 = ~n1114 & n1153;
  assign n1155 = ~n1131 & n1154;
  assign po001 = ~n1148 & n1155;
  assign n1157 = ~n695 & ~po078;
  assign n1158 = n695 & po078;
  assign n1159 = ~n1157 & ~n1158;
  assign n1160 = ~n795 & ~po080;
  assign n1161 = n795 & po080;
  assign n1162 = ~n1160 & ~n1161;
  assign n1163 = ~n863 & ~po081;
  assign n1164 = n863 & po081;
  assign n1165 = ~n1163 & ~n1164;
  assign n1166 = ~n802 & ~po079;
  assign n1167 = n802 & po079;
  assign n1168 = ~n1166 & ~n1167;
  assign n1169 = ~n673 & n1159;
  assign n1170 = n1162 & n1169;
  assign n1171 = n1165 & n1170;
  assign n1172 = n1168 & n1171;
  assign n1173 = pi083 & n1172;
  assign n1174 = ~po078 & ~n923;
  assign n1175 = po078 & n923;
  assign n1176 = ~n1174 & ~n1175;
  assign n1177 = ~po080 & ~n946;
  assign n1178 = po080 & n946;
  assign n1179 = ~n1177 & ~n1178;
  assign n1180 = ~po081 & ~n976;
  assign n1181 = po081 & n976;
  assign n1182 = ~n1180 & ~n1181;
  assign n1183 = ~po079 & ~n953;
  assign n1184 = po079 & n953;
  assign n1185 = ~n1183 & ~n1184;
  assign n1186 = ~n673 & n1176;
  assign n1187 = n1179 & n1186;
  assign n1188 = n1182 & n1187;
  assign n1189 = n1185 & n1188;
  assign n1190 = pi082 & n1189;
  assign n1191 = ~po078 & ~n1008;
  assign n1192 = po078 & n1008;
  assign n1193 = ~n1191 & ~n1192;
  assign n1194 = ~po080 & ~n1031;
  assign n1195 = po080 & n1031;
  assign n1196 = ~n1194 & ~n1195;
  assign n1197 = ~po081 & ~n1061;
  assign n1198 = po081 & n1061;
  assign n1199 = ~n1197 & ~n1198;
  assign n1200 = ~po079 & ~n1038;
  assign n1201 = po079 & n1038;
  assign n1202 = ~n1200 & ~n1201;
  assign n1203 = ~n673 & n1193;
  assign n1204 = n1196 & n1203;
  assign n1205 = n1199 & n1204;
  assign n1206 = n1202 & n1205;
  assign n1207 = pi081 & n1206;
  assign n1208 = ~n673 & po078;
  assign n1209 = ~po080 & n1208;
  assign n1210 = ~po081 & n1209;
  assign n1211 = ~po079 & n1210;
  assign n1212 = pi010 & n1211;
  assign n1213 = ~n673 & ~po080;
  assign n1214 = ~po081 & n1213;
  assign n1215 = po079 & n1214;
  assign n1216 = po078 & n1215;
  assign n1217 = pi010 & n1216;
  assign n1218 = pi011 & n1217;
  assign n1219 = ~n681 & ~po078;
  assign n1220 = n681 & po078;
  assign n1221 = ~n1219 & ~n1220;
  assign n1222 = ~n760 & ~po080;
  assign n1223 = n760 & po080;
  assign n1224 = ~n1222 & ~n1223;
  assign n1225 = ~n834 & ~po081;
  assign n1226 = n834 & po081;
  assign n1227 = ~n1225 & ~n1226;
  assign n1228 = ~n727 & ~po079;
  assign n1229 = n727 & po079;
  assign n1230 = ~n1228 & ~n1229;
  assign n1231 = ~n673 & n1221;
  assign n1232 = n1224 & n1231;
  assign n1233 = n1227 & n1232;
  assign n1234 = n1230 & n1233;
  assign n1235 = n753 & n1234;
  assign n1236 = ~n684 & ~po078;
  assign n1237 = n684 & po078;
  assign n1238 = ~n1236 & ~n1237;
  assign n1239 = ~n766 & ~po080;
  assign n1240 = n766 & po080;
  assign n1241 = ~n1239 & ~n1240;
  assign n1242 = ~n842 & ~po081;
  assign n1243 = n842 & po081;
  assign n1244 = ~n1242 & ~n1243;
  assign n1245 = ~n734 & ~po079;
  assign n1246 = n734 & po079;
  assign n1247 = ~n1245 & ~n1246;
  assign n1248 = ~n673 & n1238;
  assign n1249 = n1241 & n1248;
  assign n1250 = n1244 & n1249;
  assign n1251 = n1247 & n1250;
  assign n1252 = n747 & n1251;
  assign n1253 = ~n687 & ~po078;
  assign n1254 = n687 & po078;
  assign n1255 = ~n1253 & ~n1254;
  assign n1256 = ~n772 & ~po080;
  assign n1257 = n772 & po080;
  assign n1258 = ~n1256 & ~n1257;
  assign n1259 = ~n850 & ~po081;
  assign n1260 = n850 & po081;
  assign n1261 = ~n1259 & ~n1260;
  assign n1262 = ~n782 & ~po079;
  assign n1263 = n782 & po079;
  assign n1264 = ~n1262 & ~n1263;
  assign n1265 = ~n673 & n1255;
  assign n1266 = n1258 & n1265;
  assign n1267 = n1261 & n1266;
  assign n1268 = n1264 & n1267;
  assign n1269 = n741 & n1268;
  assign n1270 = n534 & ~n1173;
  assign n1271 = ~n1190 & n1270;
  assign n1272 = ~n1207 & n1271;
  assign n1273 = ~n1212 & n1272;
  assign n1274 = ~n1218 & n1273;
  assign n1275 = ~n1235 & n1274;
  assign n1276 = ~n1252 & n1275;
  assign po002 = ~n1269 & n1276;
  assign po003 = pi006 & pi007;
  assign n1279 = pi043 & pi181;
  assign n1280 = ~pi007 & n1279;
  assign n1281 = pi052 & ~n1280;
  assign po062 = pi074 & n1281;
  assign po099 = pi052 & pi074;
  assign po095 = pi052 & pi149;
  assign po118 = pi052 & pi162;
  assign po056 = pi052 & pi071;
  assign po054 = pi052 & pi070;
  assign po061 = pi031 & pi052;
  assign n1289 = ~pi007 & pi166;
  assign po120 = pi030 & pi052;
  assign po124 = ~n1289 & po120;
  assign po094 = pi052 & pi148;
  assign n1293 = ~po061 & ~po124;
  assign n1294 = ~po094 & n1293;
  assign n1295 = ~po120 & n1294;
  assign n1296 = ~po118 & ~po056;
  assign n1297 = ~po054 & n1296;
  assign n1298 = ~po062 & ~po099;
  assign n1299 = ~po095 & n1298;
  assign n1300 = n1297 & n1299;
  assign po004 = ~n1295 | ~n1300;
  assign n1302 = pi009 & pi064;
  assign n1303 = ~pi058 & n1302;
  assign n1304 = pi059 & n1303;
  assign n1305 = ~pi008 & ~n1304;
  assign po005 = pi009 & ~n1305;
  assign n1307 = pi033 & pi034;
  assign n1308 = pi035 & n1307;
  assign n1309 = pi036 & n1308;
  assign n1310 = pi058 & ~pi059;
  assign n1311 = pi064 & n1310;
  assign n1312 = pi199 & ~n1311;
  assign po160 = ~pi177 & n1312;
  assign n1314 = ~pi012 & n1309;
  assign n1315 = po160 & n1314;
  assign n1316 = pi037 & n1315;
  assign n1317 = n534 & ~n1091;
  assign n1318 = ~n1212 & n1317;
  assign n1319 = n534 & ~n1097;
  assign n1320 = ~n1218 & n1319;
  assign n1321 = n1318 & n1320;
  assign n1322 = pi010 & ~n1321;
  assign n1323 = pi011 & n1322;
  assign n1324 = n534 & ~n1001;
  assign n1325 = ~n1190 & n1324;
  assign n1326 = n534 & ~n1131;
  assign n1327 = ~n1252 & n1326;
  assign n1328 = n1325 & n1327;
  assign n1329 = n747 & ~n1328;
  assign n1330 = n534 & ~n916;
  assign n1331 = ~n1173 & n1330;
  assign n1332 = n534 & ~n1148;
  assign n1333 = ~n1269 & n1332;
  assign n1334 = n1331 & n1333;
  assign n1335 = n741 & ~n1334;
  assign n1336 = n534 & ~n1086;
  assign n1337 = ~n1207 & n1336;
  assign n1338 = n534 & ~n1114;
  assign n1339 = ~n1235 & n1338;
  assign n1340 = n1337 & n1339;
  assign n1341 = n753 & ~n1340;
  assign n1342 = ~n1335 & ~n1341;
  assign n1343 = ~n1323 & ~n1329;
  assign n1344 = n1342 & n1343;
  assign n1345 = pi110 & ~n545;
  assign n1346 = n567 & n1345;
  assign n1347 = pi120 & n545;
  assign n1348 = ~n567 & n1347;
  assign n1349 = ~n1346 & ~n1348;
  assign n1350 = ~n557 & ~n1349;
  assign n1351 = n534 & n1350;
  assign n1352 = ~n542 & n1351;
  assign n1353 = ~n578 & n1352;
  assign n1354 = ~n578 & n1353;
  assign n1355 = pi136 & n583;
  assign n1356 = n578 & n1355;
  assign n1357 = n578 & n1356;
  assign n1358 = ~n1354 & ~n1357;
  assign n1359 = ~n662 & ~n1358;
  assign n1360 = n661 & n1359;
  assign n1361 = pi139 & n662;
  assign n1362 = ~n661 & n1361;
  assign po083 = n1360 | n1362;
  assign n1364 = pi111 & ~n545;
  assign n1365 = n567 & n1364;
  assign n1366 = pi121 & n545;
  assign n1367 = ~n567 & n1366;
  assign n1368 = ~n1365 & ~n1367;
  assign n1369 = ~n557 & ~n1368;
  assign n1370 = n534 & n1369;
  assign n1371 = ~n542 & n1370;
  assign n1372 = ~n578 & n1371;
  assign n1373 = ~n578 & n1372;
  assign n1374 = pi137 & n583;
  assign n1375 = n578 & n1374;
  assign n1376 = n578 & n1375;
  assign n1377 = ~n1373 & ~n1376;
  assign n1378 = ~n662 & ~n1377;
  assign n1379 = n661 & n1378;
  assign n1380 = pi140 & n662;
  assign n1381 = ~n661 & n1380;
  assign po084 = n1379 | n1381;
  assign n1383 = pi109 & ~n545;
  assign n1384 = n567 & n1383;
  assign n1385 = pi119 & n545;
  assign n1386 = ~n567 & n1385;
  assign n1387 = ~n1384 & ~n1386;
  assign n1388 = ~n557 & ~n1387;
  assign n1389 = n534 & n1388;
  assign n1390 = ~n542 & n1389;
  assign n1391 = ~n578 & n1390;
  assign n1392 = ~n578 & n1391;
  assign n1393 = pi135 & n583;
  assign n1394 = n578 & n1393;
  assign n1395 = n578 & n1394;
  assign n1396 = ~n1392 & ~n1395;
  assign n1397 = ~n662 & ~n1396;
  assign n1398 = n661 & n1397;
  assign n1399 = pi138 & n662;
  assign n1400 = ~n661 & n1399;
  assign po082 = n1398 | n1400;
  assign n1402 = ~pi012 & ~n1344;
  assign n1403 = po083 & n1402;
  assign n1404 = po084 & n1403;
  assign n1405 = po082 & n1404;
  assign n1406 = po160 & n1405;
  assign n1407 = pi119 & pi121;
  assign n1408 = pi123 & n1407;
  assign n1409 = pi125 & n1408;
  assign n1410 = pi127 & n1409;
  assign n1411 = pi126 & n1410;
  assign n1412 = pi124 & n1411;
  assign n1413 = pi122 & n1412;
  assign n1414 = pi120 & n1413;
  assign n1415 = ~pi012 & n1414;
  assign n1416 = po160 & n1415;
  assign n1417 = ~n1316 & ~n1406;
  assign po006 = n1416 | ~n1417;
  assign n1419 = ~po052 & ~n627;
  assign n1420 = po065 & ~n1419;
  assign n1421 = ~n540 & ~n567;
  assign n1422 = po065 & n1421;
  assign n1423 = pi018 & ~n1311;
  assign n1424 = po052 & n1423;
  assign n1425 = ~pi017 & n1424;
  assign n1426 = pi029 & n644;
  assign n1427 = pi066 & n603;
  assign n1428 = ~pi066 & n616;
  assign n1429 = ~n1427 & ~n1428;
  assign n1430 = ~n627 & ~n1429;
  assign n1431 = ~n1426 & ~n1430;
  assign n1432 = ~pi016 & ~n631;
  assign n1433 = ~n628 & n1431;
  assign n1434 = n1432 & n1433;
  assign n1435 = pi004 & ~n1434;
  assign n1436 = n534 & n647;
  assign n1437 = ~n630 & n1436;
  assign n1438 = n648 & n1437;
  assign n1439 = po065 & ~n1438;
  assign n1440 = n627 & ~n1429;
  assign n1441 = ~n626 & ~n627;
  assign n1442 = n647 & ~n1440;
  assign n1443 = ~n1441 & n1442;
  assign n1444 = n534 & n1443;
  assign n1445 = pi015 & ~n1444;
  assign n1446 = pi014 & n628;
  assign n1447 = pi019 & ~n534;
  assign n1448 = ~n1425 & ~n1435;
  assign n1449 = ~po160 & ~n1422;
  assign n1450 = n1448 & n1449;
  assign n1451 = ~n1446 & ~n1447;
  assign n1452 = ~n1439 & ~n1445;
  assign n1453 = n1451 & n1452;
  assign po009 = ~n1450 | ~n1453;
  assign n1455 = pi012 & po160;
  assign n1456 = ~po009 & ~n1455;
  assign n1457 = ~pi063 & n1311;
  assign n1458 = po160 & n1457;
  assign n1459 = pi039 & po160;
  assign n1460 = n1304 & po160;
  assign n1461 = ~pi021 & ~n1420;
  assign n1462 = ~n1456 & n1461;
  assign n1463 = ~pi020 & n1462;
  assign n1464 = ~n1458 & n1463;
  assign n1465 = ~n1459 & n1464;
  assign n1466 = ~n1416 & n1465;
  assign n1467 = ~n1406 & n1466;
  assign n1468 = ~n1460 & n1467;
  assign po007 = n1316 | ~n1468;
  assign n1470 = pi004 & ~n1431;
  assign n1471 = pi015 & ~n1443;
  assign n1472 = ~n1446 & ~n1470;
  assign n1473 = ~n1471 & n1472;
  assign n1474 = ~pi203 & pi204;
  assign n1475 = pi203 & pi204;
  assign po165 = n1474 | n1475;
  assign n1477 = ~n1311 & ~n1473;
  assign po008 = po165 | ~n1477;
  assign n1479 = pi017 & pi018;
  assign n1480 = ~pi002 & ~n782;
  assign n1481 = pi002 & n782;
  assign n1482 = ~n1480 & ~n1481;
  assign n1483 = ~pi000 & ~n850;
  assign n1484 = pi000 & n850;
  assign n1485 = ~n1483 & ~n1484;
  assign n1486 = ~pi001 & ~n772;
  assign n1487 = pi001 & n772;
  assign n1488 = ~n1486 & ~n1487;
  assign n1489 = n1482 & n1485;
  assign n1490 = pi003 & n1489;
  assign n1491 = n687 & n1490;
  assign n1492 = n1488 & n1491;
  assign n1493 = pi001 & n1485;
  assign n1494 = n772 & n1493;
  assign n1495 = n782 & n1488;
  assign n1496 = pi002 & n1495;
  assign n1497 = n1485 & n1496;
  assign n1498 = ~n1484 & ~n1497;
  assign n1499 = ~n1492 & ~n1494;
  assign n1500 = n1498 & n1499;
  assign n1501 = pi018 & po052;
  assign n1502 = ~pi029 & n596;
  assign n1503 = pi027 & n1502;
  assign n1504 = pi018 & n1503;
  assign n1505 = ~n538 & ~n599;
  assign n1506 = po065 & ~n1505;
  assign n1507 = ~po052 & n1506;
  assign n1508 = po065 & n544;
  assign n1509 = ~pi016 & n494;
  assign n1510 = ~pi029 & n497;
  assign n1511 = pi027 & n1510;
  assign n1512 = ~pi029 & n492;
  assign n1513 = pi027 & n1512;
  assign n1514 = ~pi027 & n1512;
  assign n1515 = ~n1513 & ~n1514;
  assign n1516 = ~n1509 & ~n1511;
  assign n1517 = n1515 & n1516;
  assign n1518 = pi004 & ~n1517;
  assign n1519 = ~n1508 & ~n1518;
  assign n1520 = ~n1501 & ~n1504;
  assign n1521 = ~n1507 & n1520;
  assign n1522 = n1519 & n1521;
  assign n1523 = ~n1500 & ~n1522;
  assign n1524 = ~pi065 & pi066;
  assign n1525 = pi065 & ~pi066;
  assign n1526 = ~n1524 & ~n1525;
  assign n1527 = pi138 & ~pi139;
  assign n1528 = ~pi138 & pi139;
  assign n1529 = ~n1527 & ~n1528;
  assign n1530 = ~n1526 & n1529;
  assign n1531 = n1526 & ~n1529;
  assign n1532 = ~n1530 & ~n1531;
  assign n1533 = pi140 & ~pi141;
  assign n1534 = ~pi140 & pi141;
  assign n1535 = ~n1533 & ~n1534;
  assign n1536 = pi142 & ~pi143;
  assign n1537 = ~pi142 & pi143;
  assign n1538 = ~n1536 & ~n1537;
  assign n1539 = ~n1535 & n1538;
  assign n1540 = n1535 & ~n1538;
  assign n1541 = ~n1539 & ~n1540;
  assign n1542 = ~n1532 & n1541;
  assign n1543 = n1532 & ~n1541;
  assign n1544 = ~n1542 & ~n1543;
  assign n1545 = pi256 & n1544;
  assign n1546 = ~pi256 & ~n1544;
  assign n1547 = ~n1545 & ~n1546;
  assign n1548 = pi144 & ~pi145;
  assign n1549 = ~pi144 & pi145;
  assign n1550 = ~n1548 & ~n1549;
  assign n1551 = pi146 & ~pi147;
  assign n1552 = ~pi146 & pi147;
  assign n1553 = ~n1551 & ~n1552;
  assign n1554 = ~n1550 & n1553;
  assign n1555 = n1550 & ~n1553;
  assign n1556 = ~n1554 & ~n1555;
  assign n1557 = ~pi246 & pi247;
  assign n1558 = pi246 & ~pi247;
  assign n1559 = ~n1557 & ~n1558;
  assign n1560 = pi253 & ~pi254;
  assign n1561 = ~pi253 & pi254;
  assign n1562 = ~n1560 & ~n1561;
  assign n1563 = ~n1559 & n1562;
  assign n1564 = n1559 & ~n1562;
  assign n1565 = ~n1563 & ~n1564;
  assign n1566 = ~n1556 & n1565;
  assign n1567 = n1556 & ~n1565;
  assign n1568 = ~n1566 & ~n1567;
  assign n1569 = pi255 & n1568;
  assign n1570 = ~pi255 & ~n1568;
  assign n1571 = ~n1569 & ~n1570;
  assign n1572 = ~n1547 & ~n1571;
  assign n1573 = ~pi056 & n668;
  assign n1574 = n489 & n1573;
  assign n1575 = pi029 & n1574;
  assign n1576 = pi027 & n1575;
  assign n1577 = ~n598 & ~n1514;
  assign n1578 = ~n1576 & n1577;
  assign n1579 = pi004 & ~n1578;
  assign n1580 = ~n544 & ~n599;
  assign n1581 = ~n538 & n1580;
  assign n1582 = po065 & ~n1581;
  assign n1583 = ~n1579 & ~n1582;
  assign n1584 = ~n1572 & ~n1583;
  assign n1585 = pi004 & pi177;
  assign n1586 = pi187 & ~n1585;
  assign n1587 = ~pi020 & ~pi021;
  assign n1588 = n534 & n1587;
  assign n1589 = ~n1479 & n1588;
  assign n1590 = ~n1523 & n1589;
  assign n1591 = ~po165 & n1590;
  assign n1592 = ~n1420 & n1591;
  assign n1593 = ~n1584 & n1592;
  assign n1594 = ~n1586 & n1593;
  assign n1595 = po009 & n1594;
  assign n1596 = ~n1458 & n1595;
  assign n1597 = ~n1459 & n1596;
  assign n1598 = ~n1416 & n1597;
  assign n1599 = ~n1406 & n1598;
  assign n1600 = ~n1460 & n1599;
  assign po010 = ~n1316 & n1600;
  assign n1602 = pi004 & n598;
  assign n1603 = pi201 & ~n566;
  assign n1604 = ~n549 & ~n1603;
  assign n1605 = pi015 & n540;
  assign n1606 = ~n1604 & n1605;
  assign n1607 = ~n538 & ~n549;
  assign n1608 = ~n537 & n1607;
  assign n1609 = n540 & ~n1608;
  assign n1610 = po065 & n1609;
  assign n1611 = ~pi040 & ~n1610;
  assign n1612 = ~n1602 & ~n1606;
  assign n1613 = n1611 & n1612;
  assign n1614 = pi014 & n598;
  assign n1615 = ~pi039 & ~n1613;
  assign po047 = ~n1614 & n1615;
  assign po011 = po010 | po047;
  assign po012 = pi023 | ~pi150;
  assign n1619 = pi015 & n631;
  assign n1620 = n1514 & ~n1584;
  assign n1621 = ~n627 & n630;
  assign n1622 = ~n537 & ~n591;
  assign n1623 = ~n538 & ~n1620;
  assign n1624 = ~n1621 & n1623;
  assign n1625 = n1622 & n1624;
  assign n1626 = pi004 & ~n1625;
  assign n1627 = pi014 & n1513;
  assign n1628 = ~n1511 & ~n1513;
  assign n1629 = pi004 & ~n1628;
  assign n1630 = ~n1627 & ~n1629;
  assign n1631 = ~n1619 & ~n1626;
  assign po013 = ~n1630 | ~n1631;
  assign n1633 = ~pi020 & pi025;
  assign po014 = pi024 | n1633;
  assign n1635 = pi250 & ~pi251;
  assign n1636 = ~pi250 & pi251;
  assign n1637 = ~n1635 & ~n1636;
  assign n1638 = pi248 & ~pi249;
  assign n1639 = ~pi248 & pi249;
  assign n1640 = ~n1638 & ~n1639;
  assign po015 = n1637 & n1640;
  assign n1642 = pi015 & ~n627;
  assign n1643 = ~n626 & n1642;
  assign n1644 = pi004 & n1426;
  assign n1645 = pi004 & n1430;
  assign n1646 = pi015 & n1440;
  assign n1647 = pi015 & ~n647;
  assign n1648 = ~n1446 & ~n1643;
  assign n1649 = ~n1644 & n1648;
  assign n1650 = ~n1645 & n1649;
  assign n1651 = ~n1646 & n1650;
  assign n1652 = ~n1647 & n1651;
  assign n1653 = ~pi021 & ~n1586;
  assign n1654 = ~n1652 & n1653;
  assign n1655 = ~n1311 & n1654;
  assign po016 = ~pi020 & n1655;
  assign po017 = n538 & po081;
  assign po018 = n538 & po080;
  assign po019 = n538 & po079;
  assign po020 = n538 & po078;
  assign n1661 = pi051 & ~n534;
  assign n1662 = ~n542 & n1661;
  assign n1663 = n557 & n1662;
  assign n1664 = pi092 & ~n545;
  assign n1665 = n567 & n1664;
  assign n1666 = pi104 & n545;
  assign n1667 = ~n567 & n1666;
  assign n1668 = ~n1665 & ~n1667;
  assign n1669 = n534 & ~n1668;
  assign n1670 = ~n542 & n1669;
  assign n1671 = ~n557 & n1670;
  assign n1672 = ~n1663 & ~n1671;
  assign n1673 = ~n578 & ~n1672;
  assign n1674 = ~n578 & n1673;
  assign n1675 = ~n662 & n1674;
  assign n1676 = n661 & n1675;
  assign n1677 = pi134 & n662;
  assign n1678 = ~n661 & n1677;
  assign po077 = n1676 | n1678;
  assign po021 = n538 & po077;
  assign n1681 = pi129 & ~n534;
  assign n1682 = ~n542 & n1681;
  assign n1683 = n557 & n1682;
  assign n1684 = pi091 & ~n545;
  assign n1685 = n567 & n1684;
  assign n1686 = pi103 & n545;
  assign n1687 = ~n567 & n1686;
  assign n1688 = ~n1685 & ~n1687;
  assign n1689 = n534 & ~n1688;
  assign n1690 = ~n542 & n1689;
  assign n1691 = ~n557 & n1690;
  assign n1692 = ~n1683 & ~n1691;
  assign n1693 = ~n578 & ~n1692;
  assign n1694 = ~n578 & n1693;
  assign n1695 = n578 & ~n583;
  assign n1696 = n578 & n1695;
  assign n1697 = ~n1694 & ~n1696;
  assign n1698 = ~n662 & ~n1697;
  assign n1699 = n661 & n1698;
  assign n1700 = pi133 & n662;
  assign n1701 = ~n661 & n1700;
  assign po076 = n1699 | n1701;
  assign po022 = n538 & po076;
  assign n1704 = pi048 & ~n534;
  assign n1705 = ~n542 & n1704;
  assign n1706 = n557 & n1705;
  assign n1707 = pi090 & ~n545;
  assign n1708 = n567 & n1707;
  assign n1709 = pi102 & n545;
  assign n1710 = ~n567 & n1709;
  assign n1711 = ~n1708 & ~n1710;
  assign n1712 = n534 & ~n1711;
  assign n1713 = ~n542 & n1712;
  assign n1714 = ~n557 & n1713;
  assign n1715 = ~n1706 & ~n1714;
  assign n1716 = ~n578 & ~n1715;
  assign n1717 = ~n578 & n1716;
  assign n1718 = n578 & n583;
  assign n1719 = n578 & n1718;
  assign n1720 = ~n1717 & ~n1719;
  assign n1721 = ~n662 & ~n1720;
  assign n1722 = n661 & n1721;
  assign n1723 = pi132 & n662;
  assign n1724 = ~n661 & n1723;
  assign po075 = n1722 | n1724;
  assign po023 = n538 & po075;
  assign n1727 = pi049 & ~n534;
  assign n1728 = ~n542 & n1727;
  assign n1729 = n557 & n1728;
  assign n1730 = pi089 & ~n545;
  assign n1731 = n567 & n1730;
  assign n1732 = pi101 & n545;
  assign n1733 = ~n567 & n1732;
  assign n1734 = ~n1731 & ~n1733;
  assign n1735 = n534 & ~n1734;
  assign n1736 = ~n542 & n1735;
  assign n1737 = ~n557 & n1736;
  assign n1738 = ~n1729 & ~n1737;
  assign n1739 = ~n578 & ~n1738;
  assign n1740 = ~n578 & n1739;
  assign n1741 = pi000 & ~n583;
  assign n1742 = ~n583 & n1741;
  assign n1743 = ~n583 & ~n1742;
  assign n1744 = n578 & ~n1743;
  assign n1745 = n578 & n1744;
  assign n1746 = ~n1740 & ~n1745;
  assign n1747 = ~n662 & ~n1746;
  assign n1748 = n661 & n1747;
  assign n1749 = pi131 & n662;
  assign n1750 = ~n661 & n1749;
  assign po074 = n1748 | n1750;
  assign po024 = n538 & po074;
  assign n1753 = pi047 & ~n534;
  assign n1754 = ~n542 & n1753;
  assign n1755 = n557 & n1754;
  assign n1756 = pi088 & ~n545;
  assign n1757 = n567 & n1756;
  assign n1758 = pi100 & n545;
  assign n1759 = ~n567 & n1758;
  assign n1760 = ~n1757 & ~n1759;
  assign n1761 = n534 & ~n1760;
  assign n1762 = ~n542 & n1761;
  assign n1763 = ~n557 & n1762;
  assign n1764 = ~n1755 & ~n1763;
  assign n1765 = ~n578 & ~n1764;
  assign n1766 = ~n578 & n1765;
  assign n1767 = pi001 & ~n583;
  assign n1768 = ~n583 & n1767;
  assign n1769 = ~n583 & ~n1768;
  assign n1770 = n578 & ~n1769;
  assign n1771 = n578 & n1770;
  assign n1772 = ~n1766 & ~n1771;
  assign n1773 = ~n662 & ~n1772;
  assign n1774 = n661 & n1773;
  assign n1775 = pi130 & n662;
  assign n1776 = ~n661 & n1775;
  assign po073 = n1774 | n1776;
  assign po025 = n538 & po073;
  assign n1779 = pi050 & ~n534;
  assign n1780 = ~n542 & n1779;
  assign n1781 = n557 & n1780;
  assign n1782 = pi087 & ~n545;
  assign n1783 = n567 & n1782;
  assign n1784 = pi099 & n545;
  assign n1785 = ~n567 & n1784;
  assign n1786 = ~n1783 & ~n1785;
  assign n1787 = n534 & ~n1786;
  assign n1788 = ~n542 & n1787;
  assign n1789 = ~n557 & n1788;
  assign n1790 = ~n1781 & ~n1789;
  assign n1791 = ~n578 & ~n1790;
  assign n1792 = ~n578 & n1791;
  assign n1793 = pi002 & ~n583;
  assign n1794 = ~n583 & n1793;
  assign n1795 = ~n583 & ~n1794;
  assign n1796 = n578 & ~n1795;
  assign n1797 = n578 & n1796;
  assign n1798 = ~n1792 & ~n1797;
  assign n1799 = ~n662 & ~n1798;
  assign n1800 = n661 & n1799;
  assign n1801 = pi137 & n662;
  assign n1802 = ~n661 & n1801;
  assign po072 = n1800 | n1802;
  assign po026 = n538 & po072;
  assign n1805 = pi046 & ~n534;
  assign n1806 = ~n542 & n1805;
  assign n1807 = n557 & n1806;
  assign n1808 = pi086 & ~n545;
  assign n1809 = n567 & n1808;
  assign n1810 = pi098 & n545;
  assign n1811 = ~n567 & n1810;
  assign n1812 = ~n1809 & ~n1811;
  assign n1813 = n534 & ~n1812;
  assign n1814 = ~n542 & n1813;
  assign n1815 = ~n557 & n1814;
  assign n1816 = ~n1807 & ~n1815;
  assign n1817 = ~n578 & ~n1816;
  assign n1818 = ~n578 & n1817;
  assign n1819 = pi000 & n583;
  assign n1820 = pi003 & ~n583;
  assign n1821 = ~n583 & n1820;
  assign n1822 = ~n1819 & ~n1821;
  assign n1823 = n578 & ~n1822;
  assign n1824 = n578 & n1823;
  assign n1825 = ~n1818 & ~n1824;
  assign n1826 = ~n662 & ~n1825;
  assign n1827 = n661 & n1826;
  assign n1828 = pi136 & n662;
  assign n1829 = ~n661 & n1828;
  assign po071 = n1827 | n1829;
  assign po027 = n538 & po071;
  assign n1832 = pi085 & ~n545;
  assign n1833 = n567 & n1832;
  assign n1834 = pi097 & n545;
  assign n1835 = ~n567 & n1834;
  assign n1836 = ~n1833 & ~n1835;
  assign n1837 = n534 & ~n1836;
  assign n1838 = ~n542 & n1837;
  assign n1839 = ~n557 & n1838;
  assign n1840 = ~n1663 & ~n1839;
  assign n1841 = ~n578 & ~n1840;
  assign n1842 = ~n578 & n1841;
  assign n1843 = pi001 & n583;
  assign n1844 = pi134 & ~n583;
  assign n1845 = ~n583 & n1844;
  assign n1846 = ~n1843 & ~n1845;
  assign n1847 = n578 & ~n1846;
  assign n1848 = n578 & n1847;
  assign n1849 = ~n1842 & ~n1848;
  assign n1850 = ~n662 & ~n1849;
  assign n1851 = n661 & n1850;
  assign n1852 = pi135 & n662;
  assign n1853 = ~n661 & n1852;
  assign po070 = n1851 | n1853;
  assign po028 = n538 & po070;
  assign n1856 = ~po065 & ~n540;
  assign n1857 = ~n567 & n1856;
  assign n1858 = pi128 & n1414;
  assign n1859 = pi023 & ~n598;
  assign n1860 = ~pi042 & n1859;
  assign n1861 = ~n1858 & n1860;
  assign n1862 = n540 & n1861;
  assign n1863 = pi244 & n1862;
  assign n1864 = pi243 & n1863;
  assign n1865 = ~n1857 & ~n1864;
  assign n1866 = po065 & n537;
  assign n1867 = po065 & po082;
  assign n1868 = n538 & n1867;
  assign n1869 = n1865 & n1868;
  assign n1870 = ~n1866 & n1869;
  assign n1871 = po065 & n538;
  assign n1872 = ~pi119 & ~n1866;
  assign n1873 = ~n1865 & n1872;
  assign n1874 = ~n1871 & n1873;
  assign po029 = n1870 | n1874;
  assign n1876 = po065 & po083;
  assign n1877 = n538 & n1876;
  assign n1878 = n1865 & n1877;
  assign n1879 = ~n1866 & n1878;
  assign n1880 = ~pi119 & pi120;
  assign n1881 = pi119 & ~pi120;
  assign n1882 = ~n1880 & ~n1881;
  assign n1883 = ~n1866 & ~n1882;
  assign n1884 = ~n1865 & n1883;
  assign n1885 = ~n1871 & n1884;
  assign po030 = n1879 | n1885;
  assign n1887 = po065 & po084;
  assign n1888 = n538 & n1887;
  assign n1889 = n1865 & n1888;
  assign n1890 = ~n1866 & n1889;
  assign n1891 = pi119 & pi120;
  assign n1892 = pi121 & ~n1891;
  assign n1893 = ~pi121 & n1891;
  assign n1894 = ~n1892 & ~n1893;
  assign n1895 = ~n1866 & ~n1894;
  assign n1896 = ~n1865 & n1895;
  assign n1897 = ~n1871 & n1896;
  assign po031 = n1890 | n1897;
  assign n1899 = pi112 & ~n545;
  assign n1900 = n567 & n1899;
  assign n1901 = pi122 & n545;
  assign n1902 = ~n567 & n1901;
  assign n1903 = ~n1900 & ~n1902;
  assign n1904 = ~n557 & ~n1903;
  assign n1905 = n534 & n1904;
  assign n1906 = ~n542 & n1905;
  assign n1907 = ~n578 & n1906;
  assign n1908 = ~n578 & n1907;
  assign n1909 = pi130 & n583;
  assign n1910 = pi135 & ~n583;
  assign n1911 = ~n583 & n1910;
  assign n1912 = ~n1909 & ~n1911;
  assign n1913 = n578 & ~n1912;
  assign n1914 = n578 & n1913;
  assign n1915 = ~n1908 & ~n1914;
  assign n1916 = ~n662 & ~n1915;
  assign n1917 = n661 & n1916;
  assign n1918 = pi141 & n662;
  assign n1919 = ~n661 & n1918;
  assign po085 = n1917 | n1919;
  assign n1921 = po065 & po085;
  assign n1922 = n538 & n1921;
  assign n1923 = n1865 & n1922;
  assign n1924 = ~n1866 & n1923;
  assign n1925 = pi120 & n1407;
  assign n1926 = pi122 & ~n1925;
  assign n1927 = ~pi122 & n1925;
  assign n1928 = ~n1926 & ~n1927;
  assign n1929 = ~n1866 & ~n1928;
  assign n1930 = ~n1865 & n1929;
  assign n1931 = ~n1871 & n1930;
  assign po032 = n1924 | n1931;
  assign n1933 = pi113 & ~n545;
  assign n1934 = n567 & n1933;
  assign n1935 = pi123 & n545;
  assign n1936 = ~n567 & n1935;
  assign n1937 = ~n1934 & ~n1936;
  assign n1938 = ~n557 & ~n1937;
  assign n1939 = n534 & n1938;
  assign n1940 = ~n542 & n1939;
  assign n1941 = ~n578 & n1940;
  assign n1942 = ~n578 & n1941;
  assign n1943 = pi131 & n583;
  assign n1944 = pi136 & ~n583;
  assign n1945 = ~n583 & n1944;
  assign n1946 = ~n1943 & ~n1945;
  assign n1947 = n578 & ~n1946;
  assign n1948 = n578 & n1947;
  assign n1949 = ~n1942 & ~n1948;
  assign n1950 = ~n662 & ~n1949;
  assign n1951 = n661 & n1950;
  assign n1952 = pi142 & n662;
  assign n1953 = ~n661 & n1952;
  assign po086 = n1951 | n1953;
  assign n1955 = po065 & po086;
  assign n1956 = n538 & n1955;
  assign n1957 = n1865 & n1956;
  assign n1958 = ~n1866 & n1957;
  assign n1959 = pi122 & n1407;
  assign n1960 = pi120 & n1959;
  assign n1961 = pi123 & ~n1960;
  assign n1962 = ~pi123 & n1960;
  assign n1963 = ~n1961 & ~n1962;
  assign n1964 = ~n1866 & ~n1963;
  assign n1965 = ~n1865 & n1964;
  assign n1966 = ~n1871 & n1965;
  assign po033 = n1958 | n1966;
  assign n1968 = pi114 & ~n545;
  assign n1969 = n567 & n1968;
  assign n1970 = pi124 & n545;
  assign n1971 = ~n567 & n1970;
  assign n1972 = ~n1969 & ~n1971;
  assign n1973 = ~n557 & ~n1972;
  assign n1974 = n534 & n1973;
  assign n1975 = ~n542 & n1974;
  assign n1976 = ~n578 & n1975;
  assign n1977 = ~n578 & n1976;
  assign n1978 = pi132 & n583;
  assign n1979 = pi137 & ~n583;
  assign n1980 = ~n583 & n1979;
  assign n1981 = ~n1978 & ~n1980;
  assign n1982 = n578 & ~n1981;
  assign n1983 = n578 & n1982;
  assign n1984 = ~n1977 & ~n1983;
  assign n1985 = ~n662 & ~n1984;
  assign n1986 = n661 & n1985;
  assign n1987 = pi143 & n662;
  assign n1988 = ~n661 & n1987;
  assign po087 = n1986 | n1988;
  assign n1990 = po065 & po087;
  assign n1991 = n538 & n1990;
  assign n1992 = n1865 & n1991;
  assign n1993 = ~n1866 & n1992;
  assign n1994 = pi122 & n1408;
  assign n1995 = pi120 & n1994;
  assign n1996 = pi124 & ~n1995;
  assign n1997 = ~pi124 & n1995;
  assign n1998 = ~n1996 & ~n1997;
  assign n1999 = ~n1866 & ~n1998;
  assign n2000 = ~n1865 & n1999;
  assign n2001 = ~n1871 & n2000;
  assign po034 = n1993 | n2001;
  assign n2003 = pi026 & po065;
  assign n2004 = n537 & n2003;
  assign n2005 = n1865 & n2004;
  assign n2006 = ~n1871 & n2005;
  assign n2007 = pi124 & n1408;
  assign n2008 = pi122 & n2007;
  assign n2009 = pi120 & n2008;
  assign n2010 = pi125 & ~n2009;
  assign n2011 = ~pi125 & n2009;
  assign n2012 = ~n2010 & ~n2011;
  assign n2013 = ~n1866 & ~n2012;
  assign n2014 = ~n1865 & n2013;
  assign n2015 = ~n1871 & n2014;
  assign n2016 = pi115 & ~n545;
  assign n2017 = n567 & n2016;
  assign n2018 = pi125 & n545;
  assign n2019 = ~n567 & n2018;
  assign n2020 = ~n2017 & ~n2019;
  assign n2021 = n534 & ~n2020;
  assign n2022 = ~n542 & n2021;
  assign n2023 = ~n557 & n2022;
  assign n2024 = ~pi015 & pi026;
  assign n2025 = ~n540 & n2024;
  assign n2026 = n537 & n2025;
  assign n2027 = n534 & n2026;
  assign n2028 = n557 & n2027;
  assign n2029 = ~n2023 & ~n2028;
  assign n2030 = ~n578 & ~n2029;
  assign n2031 = ~n578 & n2030;
  assign n2032 = pi133 & n583;
  assign n2033 = pi130 & ~n583;
  assign n2034 = ~n583 & n2033;
  assign n2035 = ~n2032 & ~n2034;
  assign n2036 = n578 & ~n2035;
  assign n2037 = n578 & n2036;
  assign n2038 = ~n2031 & ~n2037;
  assign n2039 = ~n662 & ~n2038;
  assign n2040 = n661 & n2039;
  assign n2041 = pi144 & n662;
  assign n2042 = ~n661 & n2041;
  assign po088 = n2040 | n2042;
  assign n2044 = po065 & po088;
  assign n2045 = n538 & n2044;
  assign n2046 = n1865 & n2045;
  assign n2047 = ~n1866 & n2046;
  assign n2048 = ~n2006 & ~n2015;
  assign po035 = n2047 | ~n2048;
  assign n2050 = pi027 & po065;
  assign n2051 = n537 & n2050;
  assign n2052 = n1865 & n2051;
  assign n2053 = ~n1871 & n2052;
  assign n2054 = pi124 & n1409;
  assign n2055 = pi122 & n2054;
  assign n2056 = pi120 & n2055;
  assign n2057 = pi126 & ~n2056;
  assign n2058 = ~pi126 & n2056;
  assign n2059 = ~n2057 & ~n2058;
  assign n2060 = ~n1866 & ~n2059;
  assign n2061 = ~n1865 & n2060;
  assign n2062 = ~n1871 & n2061;
  assign n2063 = pi116 & ~n545;
  assign n2064 = n567 & n2063;
  assign n2065 = pi126 & n545;
  assign n2066 = ~n567 & n2065;
  assign n2067 = ~n2064 & ~n2066;
  assign n2068 = n534 & ~n2067;
  assign n2069 = ~n542 & n2068;
  assign n2070 = ~n557 & n2069;
  assign n2071 = ~pi015 & pi027;
  assign n2072 = ~n540 & n2071;
  assign n2073 = n537 & n2072;
  assign n2074 = n534 & n2073;
  assign n2075 = n557 & n2074;
  assign n2076 = ~n2070 & ~n2075;
  assign n2077 = ~n578 & ~n2076;
  assign n2078 = ~n578 & n2077;
  assign n2079 = pi134 & n583;
  assign n2080 = pi131 & ~n583;
  assign n2081 = ~n583 & n2080;
  assign n2082 = ~n2079 & ~n2081;
  assign n2083 = n578 & ~n2082;
  assign n2084 = n578 & n2083;
  assign n2085 = ~n2078 & ~n2084;
  assign n2086 = ~n662 & ~n2085;
  assign n2087 = n661 & n2086;
  assign n2088 = pi145 & n662;
  assign n2089 = ~n661 & n2088;
  assign po089 = n2087 | n2089;
  assign n2091 = po065 & po089;
  assign n2092 = n538 & n2091;
  assign n2093 = n1865 & n2092;
  assign n2094 = ~n1866 & n2093;
  assign n2095 = ~n2053 & ~n2062;
  assign po036 = n2094 | ~n2095;
  assign n2097 = pi028 & po065;
  assign n2098 = n537 & n2097;
  assign n2099 = n1865 & n2098;
  assign n2100 = ~n1871 & n2099;
  assign n2101 = pi126 & n1409;
  assign n2102 = pi124 & n2101;
  assign n2103 = pi122 & n2102;
  assign n2104 = pi120 & n2103;
  assign n2105 = pi127 & ~n2104;
  assign n2106 = ~pi127 & n2104;
  assign n2107 = ~n2105 & ~n2106;
  assign n2108 = ~n1866 & ~n2107;
  assign n2109 = ~n1865 & n2108;
  assign n2110 = ~n1871 & n2109;
  assign n2111 = pi117 & ~n545;
  assign n2112 = n567 & n2111;
  assign n2113 = pi127 & n545;
  assign n2114 = ~n567 & n2113;
  assign n2115 = ~n2112 & ~n2114;
  assign n2116 = n534 & ~n2115;
  assign n2117 = ~n542 & n2116;
  assign n2118 = ~n557 & n2117;
  assign n2119 = ~pi015 & pi028;
  assign n2120 = ~n540 & n2119;
  assign n2121 = n537 & n2120;
  assign n2122 = n534 & n2121;
  assign n2123 = n557 & n2122;
  assign n2124 = ~n2118 & ~n2123;
  assign n2125 = ~n578 & ~n2124;
  assign n2126 = ~n578 & n2125;
  assign n2127 = pi003 & n583;
  assign n2128 = pi132 & ~n583;
  assign n2129 = ~n583 & n2128;
  assign n2130 = ~n2127 & ~n2129;
  assign n2131 = n578 & ~n2130;
  assign n2132 = n578 & n2131;
  assign n2133 = ~n2126 & ~n2132;
  assign n2134 = ~n662 & ~n2133;
  assign n2135 = n661 & n2134;
  assign n2136 = pi146 & n662;
  assign n2137 = ~n661 & n2136;
  assign po090 = n2135 | n2137;
  assign n2139 = po065 & po090;
  assign n2140 = n538 & n2139;
  assign n2141 = n1865 & n2140;
  assign n2142 = ~n1866 & n2141;
  assign n2143 = ~n2100 & ~n2110;
  assign po037 = n2142 | ~n2143;
  assign n2145 = pi029 & po065;
  assign n2146 = n537 & n2145;
  assign n2147 = n1865 & n2146;
  assign n2148 = ~n1871 & n2147;
  assign n2149 = pi128 & ~n1414;
  assign n2150 = ~pi128 & n1414;
  assign n2151 = ~n2149 & ~n2150;
  assign n2152 = ~n1866 & ~n2151;
  assign n2153 = ~n1865 & n2152;
  assign n2154 = ~n1871 & n2153;
  assign n2155 = po065 & ~po000;
  assign n2156 = n538 & n2155;
  assign n2157 = n1865 & n2156;
  assign n2158 = ~n1866 & n2157;
  assign n2159 = ~n2148 & ~n2154;
  assign po038 = n2158 | ~n2159;
  assign n2161 = po065 & ~n567;
  assign po040 = ~pi033 & ~n2161;
  assign n2163 = ~pi033 & pi034;
  assign n2164 = ~n2161 & n2163;
  assign n2165 = pi033 & ~pi034;
  assign n2166 = ~n2161 & n2165;
  assign po041 = n2164 | n2166;
  assign n2168 = pi035 & ~n1307;
  assign n2169 = ~n2161 & n2168;
  assign n2170 = ~pi035 & n1307;
  assign n2171 = ~n2161 & n2170;
  assign po042 = n2169 | n2171;
  assign n2173 = pi036 & ~n1308;
  assign n2174 = ~n2161 & n2173;
  assign n2175 = ~pi036 & n1308;
  assign n2176 = ~n2161 & n2175;
  assign po043 = n2174 | n2176;
  assign n2178 = pi037 & ~n1309;
  assign n2179 = ~n2161 & n2178;
  assign n2180 = ~pi037 & n1309;
  assign n2181 = ~n2161 & n2180;
  assign po044 = n2179 | n2181;
  assign n2183 = pi014 & ~pi021;
  assign n2184 = n1513 & n2183;
  assign n2185 = ~n1311 & n2184;
  assign n2186 = ~n1311 & ~n1586;
  assign n2187 = n1626 & n2186;
  assign n2188 = ~pi021 & n2187;
  assign n2189 = ~n631 & ~n1620;
  assign n2190 = pi015 & ~pi021;
  assign n2191 = ~n2189 & n2190;
  assign n2192 = ~n1311 & n2191;
  assign n2193 = ~n2185 & ~n2188;
  assign po045 = ~n2192 & n2193;
  assign n2195 = ~pi025 & pi252;
  assign n2196 = pi025 & ~pi252;
  assign n2197 = ~n2195 & ~n2196;
  assign po046 = pi038 & n2197;
  assign n2199 = pi042 & ~pi043;
  assign n2200 = ~pi023 & n2199;
  assign po049 = pi023 | n2200;
  assign n2202 = pi042 & ~po049;
  assign n2203 = pi023 & ~n2200;
  assign n2204 = pi041 & n2203;
  assign po048 = ~n2202 & ~n2204;
  assign n2206 = ~pi078 & n1311;
  assign n2207 = pi063 & n2206;
  assign n2208 = pi191 & ~n1604;
  assign n2209 = ~po065 & n2208;
  assign n2210 = pi245 & n2209;
  assign n2211 = ~pi044 & n2210;
  assign n2212 = n540 & n2211;
  assign n2213 = ~pi027 & n1510;
  assign n2214 = ~n544 & n2213;
  assign n2215 = n1586 & n2214;
  assign n2216 = pi014 & n2215;
  assign n2217 = ~n544 & n627;
  assign n2218 = n1586 & n2217;
  assign n2219 = pi015 & n2218;
  assign n2220 = pi171 & pi177;
  assign n2221 = pi017 & n2220;
  assign n2222 = ~n544 & n1586;
  assign n2223 = ~n1509 & n2222;
  assign n2224 = ~n2213 & n2223;
  assign n2225 = ~n627 & n2224;
  assign n2226 = pi015 & ~n544;
  assign n2227 = n1586 & n2226;
  assign n2228 = n1509 & n2227;
  assign n2229 = ~n2221 & ~n2225;
  assign n2230 = ~n2228 & n2229;
  assign n2231 = ~n2216 & ~n2219;
  assign n2232 = ~pi021 & n2231;
  assign n2233 = n2230 & n2232;
  assign n2234 = pi004 & ~n566;
  assign n2235 = ~n540 & ~n2234;
  assign n2236 = pi200 & n2235;
  assign n2237 = ~po065 & n2236;
  assign n2238 = ~n567 & n2237;
  assign n2239 = pi191 & ~n540;
  assign n2240 = ~n1604 & n2239;
  assign n2241 = ~po065 & n2240;
  assign n2242 = pi243 & pi244;
  assign n2243 = pi200 & n2242;
  assign n2244 = ~po065 & n2243;
  assign n2245 = pi245 & n2244;
  assign n2246 = ~pi044 & n2245;
  assign n2247 = n540 & n2246;
  assign n2248 = ~n2241 & ~n2247;
  assign n2249 = ~n2212 & n2233;
  assign n2250 = ~n2238 & n2249;
  assign n2251 = n2248 & n2250;
  assign n2252 = ~n1457 & n2251;
  assign n2253 = ~pi039 & ~n2207;
  assign n2254 = n2252 & n2253;
  assign n2255 = pi019 & ~n533;
  assign n2256 = po052 & n2255;
  assign n2257 = n2254 & n2256;
  assign po053 = pi150 & n2257;
  assign n2259 = pi006 & ~pi007;
  assign po055 = pi071 & n2259;
  assign n2261 = pi004 & ~n500;
  assign n2262 = ~pi016 & n2261;
  assign n2263 = ~pi069 & ~n2262;
  assign n2264 = pi072 & ~n2263;
  assign po057 = pi071 & n2264;
  assign po058 = pi031 & n2259;
  assign po059 = pi070 & pi073;
  assign po060 = pi031 & pi073;
  assign n2269 = ~pi026 & ~pi056;
  assign n2270 = pi029 & n2269;
  assign n2271 = n489 & n2270;
  assign n2272 = pi028 & n2271;
  assign n2273 = ~pi027 & n2272;
  assign n2274 = pi056 & n594;
  assign n2275 = n489 & n2274;
  assign n2276 = ~pi029 & n2275;
  assign n2277 = ~pi027 & n2276;
  assign n2278 = pi027 & n671;
  assign n2279 = ~n672 & ~n2277;
  assign n2280 = n489 & n2279;
  assign n2281 = pi056 & n2280;
  assign n2282 = ~n2278 & n2281;
  assign n2283 = ~pi029 & n1574;
  assign n2284 = ~pi027 & n2283;
  assign n2285 = ~n2273 & ~n2282;
  assign n2286 = ~n2284 & n2285;
  assign n2287 = ~pi039 & ~n2286;
  assign n2288 = pi053 & pi055;
  assign n2289 = pi054 & n2288;
  assign n2290 = pi053 & ~pi054;
  assign n2291 = pi055 & n2290;
  assign n2292 = pi053 & ~pi055;
  assign n2293 = pi054 & n2292;
  assign n2294 = ~n2289 & ~n2291;
  assign n2295 = n2286 & n2294;
  assign n2296 = ~n2293 & n2295;
  assign n2297 = n534 & ~n2287;
  assign n2298 = ~n2296 & n2297;
  assign n2299 = pi078 & ~n1311;
  assign n2300 = ~pi027 & n493;
  assign n2301 = ~pi027 & n1575;
  assign n2302 = ~pi015 & ~n534;
  assign n2303 = ~pi169 & n2302;
  assign n2304 = ~pi170 & n2303;
  assign n2305 = pi084 & n2304;
  assign n2306 = pi027 & n2283;
  assign n2307 = ~pi027 & n597;
  assign n2308 = ~pi027 & n1502;
  assign n2309 = ~n1576 & ~n2300;
  assign n2310 = ~n2301 & n2309;
  assign n2311 = ~n2305 & n2310;
  assign n2312 = ~n2306 & n2311;
  assign n2313 = ~n2307 & n2312;
  assign n2314 = ~n2308 & n2313;
  assign n2315 = pi004 & ~n2314;
  assign n2316 = pi077 & n1513;
  assign n2317 = ~n1511 & ~n1514;
  assign n2318 = pi014 & ~n2317;
  assign n2319 = ~n2315 & ~n2316;
  assign n2320 = ~n2318 & n2319;
  assign n2321 = ~n1311 & n2219;
  assign n2322 = pi078 & n1311;
  assign n2323 = ~n1311 & n2225;
  assign n2324 = ~n1311 & n2228;
  assign n2325 = ~n2323 & ~n2324;
  assign n2326 = ~n2216 & ~n2321;
  assign n2327 = ~n2322 & n2326;
  assign po163 = ~n2325 | ~n2327;
  assign n2329 = ~n1457 & ~n2320;
  assign n2330 = ~po163 & n2329;
  assign n2331 = ~n1304 & n2254;
  assign n2332 = ~n1604 & ~n2331;
  assign n2333 = ~pi005 & ~n2330;
  assign n2334 = ~pi039 & ~n2299;
  assign n2335 = n2333 & n2334;
  assign n2336 = ~pi021 & ~n2332;
  assign n2337 = ~n2207 & n2336;
  assign n2338 = n2335 & n2337;
  assign n2339 = pi150 & ~n2298;
  assign po063 = ~n2338 | ~n2339;
  assign po064 = n500 & n509;
  assign n2342 = po065 & n591;
  assign n2343 = ~pi079 & ~n2342;
  assign n2344 = pi028 & n2342;
  assign po066 = n2343 | n2344;
  assign n2346 = pi080 & ~n2342;
  assign n2347 = pi079 & n2346;
  assign n2348 = pi029 & n2342;
  assign n2349 = ~pi080 & n2343;
  assign n2350 = ~n2347 & ~n2348;
  assign po067 = n2349 | ~n2350;
  assign n2352 = ~n500 & n509;
  assign n2353 = pi004 & po052;
  assign n2354 = ~n500 & n2353;
  assign n2355 = ~n2263 & n2354;
  assign n2356 = po065 & ~n2298;
  assign n2357 = pi004 & ~n2286;
  assign n2358 = ~n2356 & ~n2357;
  assign n2359 = ~n2352 & ~n2355;
  assign n2360 = n2358 & n2359;
  assign n2361 = n2254 & ~n2360;
  assign po068 = pi150 & n2361;
  assign n2363 = pi014 & ~n534;
  assign n2364 = pi004 & n2286;
  assign n2365 = n2314 & n2364;
  assign n2366 = ~n2355 & n2365;
  assign n2367 = n567 & ~n591;
  assign n2368 = ~n1621 & n2367;
  assign n2369 = pi015 & ~n2368;
  assign n2370 = ~n2363 & ~n2366;
  assign n2371 = ~n2369 & n2370;
  assign n2372 = n2254 & ~n2371;
  assign po069 = pi150 & n2372;
  assign po092 = pi148 & n2259;
  assign n2375 = ~pi165 & n1514;
  assign n2376 = ~n630 & n647;
  assign n2377 = ~n538 & n2376;
  assign n2378 = ~n591 & n1429;
  assign n2379 = n626 & n2378;
  assign n2380 = n2377 & n2379;
  assign n2381 = pi165 & ~n2380;
  assign n2382 = ~pi163 & ~pi180;
  assign n2383 = n598 & ~n2382;
  assign n2384 = pi072 & pi148;
  assign n2385 = ~pi016 & n2384;
  assign n2386 = ~n2375 & n2385;
  assign n2387 = ~n2381 & n2386;
  assign n2388 = ~n2383 & n2387;
  assign po093 = ~pi008 & n2388;
  assign po096 = pi073 & pi149;
  assign po097 = ~pi014 & po096;
  assign po098 = pi074 & n2259;
  assign po100 = pi072 & pi074;
  assign po101 = pi069 & po100;
  assign po102 = pi073 & pi074;
  assign po103 = pi073 & pi148;
  assign n2397 = pi150 & n2254;
  assign n2398 = n631 & n2397;
  assign n2399 = pi014 & n2398;
  assign n2400 = ~n538 & ~n1621;
  assign n2401 = ~n537 & ~n1426;
  assign n2402 = n2400 & n2401;
  assign n2403 = ~n549 & ~n1430;
  assign n2404 = ~n591 & n2403;
  assign n2405 = n2402 & n2404;
  assign n2406 = ~pi016 & n499;
  assign n2407 = pi015 & ~po160;
  assign n2408 = ~n1509 & n2407;
  assign n2409 = n2405 & n2408;
  assign n2410 = ~n2406 & n2409;
  assign n2411 = ~n672 & n2410;
  assign n2412 = n2254 & n2411;
  assign n2413 = pi150 & n2412;
  assign po104 = n2399 | n2413;
  assign n2415 = pi004 & n2308;
  assign n2416 = ~pi039 & n544;
  assign n2417 = n599 & n627;
  assign n2418 = ~n2213 & ~n2417;
  assign n2419 = ~n1509 & ~n2416;
  assign n2420 = n2418 & n2419;
  assign n2421 = ~pi005 & pi150;
  assign n2422 = ~n2420 & n2421;
  assign n2423 = n1586 & n2422;
  assign n2424 = ~n1311 & n2423;
  assign n2425 = n485 & ~n1311;
  assign n2426 = n1586 & n2425;
  assign n2427 = ~n2424 & n2426;
  assign n2428 = ~n499 & n2427;
  assign n2429 = n485 & n2322;
  assign n2430 = ~n2428 & ~n2429;
  assign n2431 = pi150 & ~n2415;
  assign n2432 = pi151 & n2431;
  assign n2433 = n2430 & n2432;
  assign n2434 = n2430 & n2433;
  assign n2435 = ~pi061 & ~pi063;
  assign n2436 = ~pi075 & n2435;
  assign n2437 = ~pi060 & n2436;
  assign n2438 = ~pi062 & n2437;
  assign n2439 = ~n1586 & ~n2438;
  assign n2440 = ~n2430 & ~n2439;
  assign n2441 = ~n2430 & n2440;
  assign po105 = n2434 | n2441;
  assign n2443 = pi152 & n2431;
  assign n2444 = ~n2429 & n2443;
  assign n2445 = ~n2429 & n2444;
  assign n2446 = pi063 & n2429;
  assign n2447 = n2429 & n2446;
  assign po106 = n2445 | n2447;
  assign n2449 = pi153 & n2431;
  assign n2450 = ~n2429 & n2449;
  assign n2451 = ~n2429 & n2450;
  assign n2452 = pi062 & n2429;
  assign n2453 = n2429 & n2452;
  assign po107 = n2451 | n2453;
  assign n2455 = pi154 & n2431;
  assign n2456 = ~n2429 & n2455;
  assign n2457 = ~n2429 & n2456;
  assign n2458 = pi061 & n2429;
  assign n2459 = n2429 & n2458;
  assign po108 = n2457 | n2459;
  assign n2461 = pi155 & n2431;
  assign n2462 = ~n2429 & n2461;
  assign n2463 = ~n2429 & n2462;
  assign n2464 = pi060 & n2429;
  assign n2465 = n2429 & n2464;
  assign po109 = n2463 | n2465;
  assign n2467 = pi156 & n2431;
  assign n2468 = ~n2429 & n2467;
  assign n2469 = ~n2429 & n2468;
  assign n2470 = pi075 & n2429;
  assign n2471 = n2429 & n2470;
  assign po110 = n2469 | n2471;
  assign n2473 = ~n1514 & n2397;
  assign n2474 = ~n2213 & n2473;
  assign n2475 = ~n1440 & n2474;
  assign n2476 = n534 & n2475;
  assign n2477 = ~n1441 & n2476;
  assign n2478 = n647 & n2477;
  assign n2479 = ~n1511 & n2478;
  assign po111 = pi014 & n2479;
  assign n2481 = po065 & ~n566;
  assign po113 = po058 & n2481;
  assign n2483 = ~po065 & n1858;
  assign n2484 = ~po065 & n540;
  assign n2485 = pi012 & ~po065;
  assign n2486 = ~n2241 & ~n2483;
  assign n2487 = ~n566 & n2486;
  assign n2488 = ~n2484 & n2487;
  assign n2489 = ~n2485 & n2488;
  assign n2490 = ~n2241 & ~n2485;
  assign n2491 = ~n540 & n2490;
  assign n2492 = ~po065 & n2491;
  assign n2493 = n549 & n2492;
  assign n2494 = ~n1858 & n2493;
  assign n2495 = ~n1864 & ~n2489;
  assign n2496 = ~n2494 & n2495;
  assign po114 = po058 & ~n2496;
  assign n2498 = po065 & ~n1580;
  assign n2499 = ~n591 & ~n2498;
  assign n2500 = pi031 & ~n2499;
  assign po115 = n2259 & n2500;
  assign n2502 = pi004 & ~n1311;
  assign n2503 = n1576 & n2502;
  assign n2504 = ~n1584 & n2503;
  assign n2505 = pi031 & n2504;
  assign po116 = n2259 & n2505;
  assign n2507 = ~pi004 & ~pi179;
  assign n2508 = ~pi014 & n2507;
  assign n2509 = ~n534 & ~n2508;
  assign n2510 = pi031 & n2509;
  assign po117 = n2259 & n2510;
  assign n2512 = po052 & n2397;
  assign n2513 = ~pi061 & n2512;
  assign n2514 = pi075 & n2513;
  assign n2515 = ~pi060 & n2514;
  assign n2516 = pi062 & n2515;
  assign n2517 = pi019 & n2516;
  assign n2518 = ~n1513 & n2397;
  assign n2519 = pi077 & n2518;
  assign n2520 = ~n628 & n2519;
  assign po119 = n2517 | n2520;
  assign po121 = pi030 & n2259;
  assign po122 = pi030 & pi073;
  assign po123 = pi030 & pi072;
  assign n2525 = pi018 & n2254;
  assign po125 = pi150 & n2525;
  assign n2527 = pi167 & ~n538;
  assign n2528 = pi150 & n2527;
  assign po126 = n2300 | n2528;
  assign po127 = ~pi150 | n540;
  assign n2531 = pi157 & pi158;
  assign n2532 = pi159 & n2531;
  assign n2533 = pi160 & n2532;
  assign n2534 = pi161 & n2533;
  assign n2535 = pi206 & n2534;
  assign n2536 = ~n2509 & ~n2535;
  assign n2537 = pi150 & n2536;
  assign n2538 = pi084 & n2537;
  assign n2539 = pi150 & ~n2536;
  assign n2540 = ~pi084 & n2539;
  assign po128 = n2538 | n2540;
  assign n2542 = ~pi084 & n2509;
  assign n2543 = pi084 & n2535;
  assign n2544 = ~n2542 & ~n2543;
  assign n2545 = pi169 & n2544;
  assign n2546 = pi150 & n2545;
  assign n2547 = ~pi169 & ~n2544;
  assign n2548 = pi150 & n2547;
  assign po129 = n2546 | n2548;
  assign n2550 = ~pi169 & n2542;
  assign n2551 = pi169 & n2543;
  assign n2552 = ~n2550 & ~n2551;
  assign n2553 = pi170 & n2552;
  assign n2554 = pi150 & n2553;
  assign n2555 = ~pi170 & ~n2552;
  assign n2556 = pi150 & n2555;
  assign po130 = n2554 | n2556;
  assign n2558 = pi150 & ~n1503;
  assign n2559 = n2254 & n2558;
  assign po131 = pi171 & n2559;
  assign n2561 = po065 & po165;
  assign n2562 = n544 & n2561;
  assign n2563 = ~n544 & po165;
  assign n2564 = ~n1584 & ~n2562;
  assign po132 = n2563 | ~n2564;
  assign n2566 = ~pi021 & pi174;
  assign n2567 = ~pi019 & ~pi172;
  assign n2568 = ~pi018 & n2567;
  assign n2569 = ~pi173 & n2568;
  assign n2570 = pi017 & pi150;
  assign n2571 = ~n2569 & n2570;
  assign n2572 = n2233 & n2571;
  assign po134 = n2566 | n2572;
  assign n2574 = pi004 & ~n545;
  assign n2575 = pi178 & n2574;
  assign n2576 = pi168 & ~n567;
  assign n2577 = ~n2575 & ~n2576;
  assign n2578 = pi176 & n2577;
  assign n2579 = ~pi012 & n2578;
  assign n2580 = ~n1585 & n2579;
  assign n2581 = ~pi023 & ~pi042;
  assign n2582 = ~pi177 & n1470;
  assign n2583 = ~n1646 & ~n2580;
  assign n2584 = ~n2581 & n2583;
  assign n2585 = ~n2582 & n2584;
  assign n2586 = n544 & n1586;
  assign n2587 = pi004 & n544;
  assign n2588 = pi026 & n2587;
  assign n2589 = ~n2586 & ~n2588;
  assign n2590 = n2251 & ~n2585;
  assign po139 = ~n2589 | ~n2590;
  assign n2592 = n2251 & po139;
  assign n2593 = ~n1252 & ~n1269;
  assign n2594 = ~n1235 & n2593;
  assign n2595 = ~n1218 & n2594;
  assign n2596 = ~n1097 & n2595;
  assign n2597 = ~n1114 & n2596;
  assign n2598 = ~n1131 & n2597;
  assign n2599 = ~n1148 & n2598;
  assign n2600 = ~po139 & ~n2599;
  assign po136 = n2592 | n2600;
  assign n2602 = n2251 & ~n2261;
  assign n2603 = ~n2589 & n2602;
  assign n2604 = po139 & ~n2603;
  assign n2605 = ~n1173 & ~n1269;
  assign n2606 = ~n1235 & n2605;
  assign n2607 = ~n1207 & n2606;
  assign n2608 = ~n1086 & n2607;
  assign n2609 = ~n1114 & n2608;
  assign n2610 = ~n916 & n2609;
  assign n2611 = ~n1148 & n2610;
  assign n2612 = ~po139 & ~n2611;
  assign po137 = n2604 | n2612;
  assign n2614 = n2251 & n2261;
  assign n2615 = po139 & ~n2614;
  assign n2616 = ~n1252 & n2605;
  assign n2617 = ~n1190 & n2616;
  assign n2618 = ~n1001 & n2617;
  assign n2619 = ~n1131 & n2618;
  assign n2620 = ~n916 & n2619;
  assign n2621 = ~n1148 & n2620;
  assign n2622 = ~po139 & ~n2621;
  assign po138 = n2615 | n2622;
  assign n2624 = pi172 & n2254;
  assign po140 = pi150 & n2624;
  assign n2626 = ~pi173 & ~pi179;
  assign n2627 = n2254 & ~n2626;
  assign po141 = pi150 & n2627;
  assign n2629 = ~pi109 & ~po065;
  assign n2630 = n591 & n2629;
  assign n2631 = ~n2498 & n2630;
  assign n2632 = ~po065 & n591;
  assign n2633 = po082 & ~n2632;
  assign n2634 = n2498 & n2633;
  assign po142 = n2631 | n2634;
  assign n2636 = pi109 & ~pi110;
  assign n2637 = ~pi109 & pi110;
  assign n2638 = ~n2636 & ~n2637;
  assign n2639 = ~po065 & ~n2638;
  assign n2640 = n591 & n2639;
  assign n2641 = ~n2498 & n2640;
  assign n2642 = po083 & ~n2632;
  assign n2643 = n2498 & n2642;
  assign po143 = n2641 | n2643;
  assign n2645 = pi229 & n2301;
  assign n2646 = ~n2307 & n2645;
  assign po199 = ~n2278 & n2646;
  assign n2648 = pi230 & n2301;
  assign n2649 = ~n2307 & n2648;
  assign n2650 = ~n2278 & n2649;
  assign n2651 = pi216 & ~n2301;
  assign n2652 = ~n2307 & n2651;
  assign n2653 = n2278 & n2652;
  assign po206 = n2650 | n2653;
  assign n2655 = po199 & ~po206;
  assign n2656 = ~po199 & po206;
  assign n2657 = ~n2655 & ~n2656;
  assign n2658 = pi194 & n2306;
  assign n2659 = ~n2308 & n2658;
  assign n2660 = ~n2301 & n2659;
  assign n2661 = ~n2277 & n2660;
  assign n2662 = pi152 & ~n2306;
  assign n2663 = n2308 & n2662;
  assign n2664 = ~n2301 & n2663;
  assign n2665 = ~n2277 & n2664;
  assign n2666 = pi217 & ~n2306;
  assign n2667 = ~n2308 & n2666;
  assign n2668 = n2301 & n2667;
  assign n2669 = ~n2277 & n2668;
  assign n2670 = ~n2661 & ~n2665;
  assign po193 = n2669 | ~n2670;
  assign n2672 = pi195 & n2306;
  assign n2673 = ~n2308 & n2672;
  assign n2674 = ~n2301 & n2673;
  assign n2675 = ~n2277 & n2674;
  assign n2676 = pi153 & ~n2306;
  assign n2677 = n2308 & n2676;
  assign n2678 = ~n2301 & n2677;
  assign n2679 = ~n2277 & n2678;
  assign n2680 = pi218 & ~n2306;
  assign n2681 = ~n2308 & n2680;
  assign n2682 = n2301 & n2681;
  assign n2683 = ~n2277 & n2682;
  assign n2684 = pi215 & ~n2306;
  assign n2685 = ~n2308 & n2684;
  assign n2686 = ~n2301 & n2685;
  assign n2687 = n2277 & n2686;
  assign n2688 = ~n2683 & ~n2687;
  assign n2689 = ~n2675 & ~n2679;
  assign po194 = ~n2688 | ~n2689;
  assign n2691 = po193 & ~po194;
  assign n2692 = ~po193 & po194;
  assign n2693 = ~n2691 & ~n2692;
  assign n2694 = ~n2657 & n2693;
  assign n2695 = n2657 & ~n2693;
  assign n2696 = ~n2694 & ~n2695;
  assign n2697 = pi196 & n2306;
  assign n2698 = ~n2308 & n2697;
  assign n2699 = ~n2301 & n2698;
  assign n2700 = ~n2277 & n2699;
  assign n2701 = pi154 & ~n2306;
  assign n2702 = n2308 & n2701;
  assign n2703 = ~n2301 & n2702;
  assign n2704 = ~n2277 & n2703;
  assign n2705 = pi219 & ~n2306;
  assign n2706 = ~n2308 & n2705;
  assign n2707 = n2301 & n2706;
  assign n2708 = ~n2277 & n2707;
  assign n2709 = pi214 & ~n2306;
  assign n2710 = ~n2308 & n2709;
  assign n2711 = ~n2301 & n2710;
  assign n2712 = n2277 & n2711;
  assign n2713 = ~n2708 & ~n2712;
  assign n2714 = ~n2700 & ~n2704;
  assign po195 = ~n2713 | ~n2714;
  assign n2716 = pi197 & n2306;
  assign n2717 = ~n2308 & n2716;
  assign n2718 = ~n2301 & n2717;
  assign n2719 = ~n2277 & n2718;
  assign n2720 = pi155 & ~n2306;
  assign n2721 = n2308 & n2720;
  assign n2722 = ~n2301 & n2721;
  assign n2723 = ~n2277 & n2722;
  assign n2724 = pi220 & ~n2306;
  assign n2725 = ~n2308 & n2724;
  assign n2726 = n2301 & n2725;
  assign n2727 = ~n2277 & n2726;
  assign n2728 = pi213 & ~n2306;
  assign n2729 = ~n2308 & n2728;
  assign n2730 = ~n2301 & n2729;
  assign n2731 = n2277 & n2730;
  assign n2732 = ~n2727 & ~n2731;
  assign n2733 = ~n2719 & ~n2723;
  assign po196 = ~n2732 | ~n2733;
  assign n2735 = po195 & ~po196;
  assign n2736 = ~po195 & po196;
  assign n2737 = ~n2735 & ~n2736;
  assign n2738 = pi198 & n2306;
  assign n2739 = ~n2308 & n2738;
  assign n2740 = ~n2301 & n2739;
  assign n2741 = ~n2277 & n2740;
  assign n2742 = pi156 & ~n2306;
  assign n2743 = n2308 & n2742;
  assign n2744 = ~n2301 & n2743;
  assign n2745 = ~n2277 & n2744;
  assign n2746 = pi221 & ~n2306;
  assign n2747 = ~n2308 & n2746;
  assign n2748 = n2301 & n2747;
  assign n2749 = ~n2277 & n2748;
  assign n2750 = pi212 & ~n2306;
  assign n2751 = ~n2308 & n2750;
  assign n2752 = ~n2301 & n2751;
  assign n2753 = n2277 & n2752;
  assign n2754 = ~n2749 & ~n2753;
  assign n2755 = ~n2741 & ~n2745;
  assign po197 = ~n2754 | ~n2755;
  assign n2757 = pi193 & n2306;
  assign n2758 = ~n2308 & n2757;
  assign n2759 = ~n2301 & n2758;
  assign n2760 = ~n2277 & n2759;
  assign n2761 = pi151 & ~n2306;
  assign n2762 = n2308 & n2761;
  assign n2763 = ~n2301 & n2762;
  assign n2764 = ~n2277 & n2763;
  assign n2765 = pi222 & ~n2306;
  assign n2766 = ~n2308 & n2765;
  assign n2767 = n2301 & n2766;
  assign n2768 = ~n2277 & n2767;
  assign n2769 = pi211 & ~n2306;
  assign n2770 = ~n2308 & n2769;
  assign n2771 = ~n2301 & n2770;
  assign n2772 = n2277 & n2771;
  assign n2773 = ~n2768 & ~n2772;
  assign n2774 = ~n2760 & ~n2764;
  assign po198 = ~n2773 | ~n2774;
  assign n2776 = po197 & ~po198;
  assign n2777 = ~po197 & po198;
  assign n2778 = ~n2776 & ~n2777;
  assign n2779 = ~n2737 & n2778;
  assign n2780 = n2737 & ~n2778;
  assign n2781 = ~n2779 & ~n2780;
  assign n2782 = ~n2696 & n2781;
  assign n2783 = n2696 & ~n2781;
  assign po144 = ~n2782 & ~n2783;
  assign n2785 = pi237 & n2307;
  assign n2786 = n1628 & n2785;
  assign n2787 = pi239 & ~n2307;
  assign n2788 = ~n1628 & n2787;
  assign po207 = n2786 | n2788;
  assign n2790 = pi238 & n2307;
  assign n2791 = n1628 & n2790;
  assign n2792 = pi240 & ~n2307;
  assign n2793 = ~n1628 & n2792;
  assign po208 = n2791 | n2793;
  assign n2795 = po207 & ~po208;
  assign n2796 = ~po207 & po208;
  assign n2797 = ~n2795 & ~n2796;
  assign n2798 = pi223 & n2301;
  assign n2799 = ~n2307 & n2798;
  assign n2800 = ~n2278 & n2799;
  assign n2801 = pi231 & ~n2301;
  assign n2802 = n2307 & n2801;
  assign n2803 = ~n2278 & n2802;
  assign po200 = n2800 | n2803;
  assign n2805 = pi224 & n2301;
  assign n2806 = ~n2307 & n2805;
  assign n2807 = ~n2278 & n2806;
  assign n2808 = pi232 & ~n2301;
  assign n2809 = n2307 & n2808;
  assign n2810 = ~n2278 & n2809;
  assign po201 = n2807 | n2810;
  assign n2812 = po200 & ~po201;
  assign n2813 = ~po200 & po201;
  assign n2814 = ~n2812 & ~n2813;
  assign n2815 = ~n2797 & n2814;
  assign n2816 = n2797 & ~n2814;
  assign n2817 = ~n2815 & ~n2816;
  assign n2818 = pi225 & n2301;
  assign n2819 = ~n2307 & n2818;
  assign n2820 = ~n2278 & n2819;
  assign n2821 = pi233 & ~n2301;
  assign n2822 = n2307 & n2821;
  assign n2823 = ~n2278 & n2822;
  assign po202 = n2820 | n2823;
  assign n2825 = pi226 & n2301;
  assign n2826 = ~n2307 & n2825;
  assign n2827 = ~n2278 & n2826;
  assign n2828 = pi234 & ~n2301;
  assign n2829 = n2307 & n2828;
  assign n2830 = ~n2278 & n2829;
  assign po203 = n2827 | n2830;
  assign n2832 = po202 & ~po203;
  assign n2833 = ~po202 & po203;
  assign n2834 = ~n2832 & ~n2833;
  assign n2835 = pi227 & n2301;
  assign n2836 = ~n2307 & n2835;
  assign n2837 = ~n2278 & n2836;
  assign n2838 = pi235 & ~n2301;
  assign n2839 = n2307 & n2838;
  assign n2840 = ~n2278 & n2839;
  assign po204 = n2837 | n2840;
  assign n2842 = pi228 & n2301;
  assign n2843 = ~n2307 & n2842;
  assign n2844 = ~n2278 & n2843;
  assign n2845 = pi236 & ~n2301;
  assign n2846 = n2307 & n2845;
  assign n2847 = ~n2278 & n2846;
  assign po205 = n2844 | n2847;
  assign n2849 = po204 & ~po205;
  assign n2850 = ~po204 & po205;
  assign n2851 = ~n2849 & ~n2850;
  assign n2852 = ~n2834 & n2851;
  assign n2853 = n2834 & ~n2851;
  assign n2854 = ~n2852 & ~n2853;
  assign n2855 = ~n2817 & n2854;
  assign n2856 = n2817 & ~n2854;
  assign po145 = ~n2855 & ~n2856;
  assign n2858 = pi016 & n1311;
  assign n2859 = ~pi039 & pi182;
  assign n2860 = pi016 & ~n2251;
  assign n2861 = ~n2859 & ~n2860;
  assign n2862 = ~n509 & ~n2858;
  assign po146 = ~n2861 | ~n2862;
  assign n2864 = pi014 & pi185;
  assign n2865 = pi015 & pi184;
  assign n2866 = ~n2864 & ~n2865;
  assign n2867 = n1514 & ~n2866;
  assign n2868 = ~pi186 & ~n1513;
  assign n2869 = ~n1620 & n2868;
  assign n2870 = n2197 & ~n2867;
  assign po147 = n2869 | ~n2870;
  assign n2872 = pi026 & n1508;
  assign n2873 = ~n2424 & ~n2872;
  assign po148 = n1523 | ~n2873;
  assign n2875 = ~pi005 & n534;
  assign n2876 = ~pi013 & n2875;
  assign n2877 = ~n1609 & n2876;
  assign n2878 = pi188 & n2877;
  assign po149 = pi078 | ~n2878;
  assign n2880 = ~pi015 & ~pi169;
  assign n2881 = ~pi170 & n2880;
  assign n2882 = pi084 & n2881;
  assign n2883 = pi150 & pi192;
  assign n2884 = ~n2882 & n2883;
  assign n2885 = pi192 & n2884;
  assign n2886 = n533 & ~n2885;
  assign n2887 = ~n2301 & ~n2308;
  assign n2888 = ~n1576 & n2886;
  assign n2889 = n2887 & n2888;
  assign n2890 = ~n2306 & ~n2307;
  assign n2891 = ~n2300 & n2890;
  assign n2892 = n2889 & n2891;
  assign n2893 = ~pi005 & n2892;
  assign n2894 = po163 & n2893;
  assign n2895 = n2317 & n2892;
  assign n2896 = n2886 & n2895;
  assign n2897 = ~n1513 & n2896;
  assign n2898 = ~pi005 & n2320;
  assign n2899 = n2251 & n2898;
  assign n2900 = ~n2897 & n2899;
  assign n2901 = ~n2207 & n2900;
  assign n2902 = ~pi005 & n1457;
  assign n2903 = ~po065 & n2902;
  assign n2904 = ~n1504 & ~n2894;
  assign n2905 = ~n2901 & n2904;
  assign po150 = ~n2903 & n2905;
  assign po152 = ~n533 | n2884;
  assign n2908 = pi004 & n2306;
  assign n2909 = ~n487 & ~n489;
  assign n2910 = n1311 & ~n2909;
  assign n2911 = pi078 & n2910;
  assign n2912 = ~n1311 & ~n2909;
  assign n2913 = n1586 & n2912;
  assign n2914 = ~n2424 & n2913;
  assign n2915 = ~n499 & n2914;
  assign n2916 = ~n2911 & ~n2915;
  assign n2917 = pi150 & ~n2908;
  assign n2918 = pi193 & n2917;
  assign n2919 = n2916 & n2918;
  assign n2920 = n2916 & n2919;
  assign n2921 = ~n2439 & ~n2916;
  assign n2922 = ~n2916 & n2921;
  assign po153 = n2920 | n2922;
  assign n2924 = pi194 & n2917;
  assign n2925 = ~n2911 & n2924;
  assign n2926 = ~n2911 & n2925;
  assign n2927 = pi063 & n2911;
  assign n2928 = n2911 & n2927;
  assign po154 = n2926 | n2928;
  assign n2930 = pi195 & n2917;
  assign n2931 = ~n2911 & n2930;
  assign n2932 = ~n2911 & n2931;
  assign n2933 = pi062 & n2911;
  assign n2934 = n2911 & n2933;
  assign po155 = n2932 | n2934;
  assign n2936 = pi196 & n2917;
  assign n2937 = ~n2911 & n2936;
  assign n2938 = ~n2911 & n2937;
  assign n2939 = pi061 & n2911;
  assign n2940 = n2911 & n2939;
  assign po156 = n2938 | n2940;
  assign n2942 = pi197 & n2917;
  assign n2943 = ~n2911 & n2942;
  assign n2944 = ~n2911 & n2943;
  assign n2945 = pi060 & n2911;
  assign n2946 = n2911 & n2945;
  assign po157 = n2944 | n2946;
  assign n2948 = pi198 & n2917;
  assign n2949 = ~n2911 & n2948;
  assign n2950 = ~n2911 & n2949;
  assign n2951 = pi075 & n2911;
  assign n2952 = n2911 & n2951;
  assign po158 = n2950 | n2952;
  assign n2954 = ~pi080 & n591;
  assign n2955 = ~n1304 & ~n1311;
  assign n2956 = n2254 & n2955;
  assign n2957 = ~n2954 & n2956;
  assign n2958 = pi199 & n2957;
  assign n2959 = ~pi177 & n2958;
  assign n2960 = ~n591 & ~n1421;
  assign n2961 = po065 & ~n2960;
  assign po159 = n2959 | n2961;
  assign n2963 = pi150 & pi200;
  assign n2964 = n566 & n2963;
  assign n2965 = ~n567 & n1858;
  assign n2966 = ~po139 & n2965;
  assign po161 = n2964 | n2966;
  assign n2968 = n1604 & n2902;
  assign n2969 = ~po065 & n2968;
  assign po162 = ~pi078 & n2969;
  assign n2971 = pi202 & ~n499;
  assign n2972 = pi005 & n2971;
  assign po164 = n485 | ~n2972;
  assign n2974 = pi203 & ~pi204;
  assign po166 = n1474 | n2974;
  assign n2976 = n485 & n2974;
  assign n2977 = n487 & n2974;
  assign n2978 = pi004 & n2278;
  assign n2979 = pi205 & ~n2978;
  assign n2980 = pi150 & n2979;
  assign n2981 = ~n2976 & ~n2977;
  assign po167 = n2980 | ~n2981;
  assign n2983 = ~pi066 & n598;
  assign n2984 = n598 & n2983;
  assign n2985 = ~pi243 & ~n598;
  assign n2986 = ~n598 & n2985;
  assign po169 = n2984 | n2986;
  assign n2988 = ~pi065 & n598;
  assign n2989 = n598 & n2988;
  assign n2990 = ~pi244 & ~n598;
  assign n2991 = ~n598 & n2990;
  assign po170 = n2989 | n2991;
  assign n2993 = ~n598 & ~po070;
  assign n2994 = ~n598 & n2993;
  assign n2995 = ~pi247 & n598;
  assign n2996 = n598 & n2995;
  assign po171 = n2994 | n2996;
  assign n2998 = ~n598 & ~po071;
  assign n2999 = ~n598 & n2998;
  assign n3000 = ~pi246 & n598;
  assign n3001 = n598 & n3000;
  assign po172 = n2999 | n3001;
  assign n3003 = pi022 & ~po082;
  assign n3004 = pi022 & n3003;
  assign n3005 = ~pi022 & po000;
  assign n3006 = ~pi022 & n3005;
  assign po173 = n3004 | n3006;
  assign n3008 = pi022 & ~po083;
  assign n3009 = pi022 & n3008;
  assign n3010 = ~pi022 & ~po070;
  assign n3011 = ~pi022 & n3010;
  assign po174 = n3009 | n3011;
  assign n3013 = pi022 & ~po084;
  assign n3014 = pi022 & n3013;
  assign n3015 = ~pi022 & ~po071;
  assign n3016 = ~pi022 & n3015;
  assign po175 = n3014 | n3016;
  assign n3018 = pi022 & ~po085;
  assign n3019 = pi022 & n3018;
  assign n3020 = ~pi022 & ~po072;
  assign n3021 = ~pi022 & n3020;
  assign po176 = n3019 | n3021;
  assign n3023 = pi022 & ~po086;
  assign n3024 = pi022 & n3023;
  assign n3025 = ~pi022 & ~po073;
  assign n3026 = ~pi022 & n3025;
  assign po177 = n3024 | n3026;
  assign n3028 = pi022 & ~po087;
  assign n3029 = pi022 & n3028;
  assign n3030 = ~pi022 & ~po074;
  assign n3031 = ~pi022 & n3030;
  assign po178 = n3029 | n3031;
  assign n3033 = pi022 & ~po088;
  assign n3034 = pi022 & n3033;
  assign n3035 = ~pi022 & ~po075;
  assign n3036 = ~pi022 & n3035;
  assign po179 = n3034 | n3036;
  assign n3038 = pi022 & ~po089;
  assign n3039 = pi022 & n3038;
  assign n3040 = ~pi022 & ~po076;
  assign n3041 = ~pi022 & n3040;
  assign po180 = n3039 | n3041;
  assign n3043 = pi022 & ~po090;
  assign n3044 = pi022 & n3043;
  assign n3045 = ~pi022 & ~po077;
  assign n3046 = ~pi022 & n3045;
  assign po181 = n3044 | n3046;
  assign n3048 = pi022 & ~po079;
  assign n3049 = pi022 & n3048;
  assign po182 = n3006 | n3049;
  assign n3051 = pi192 & ~n2884;
  assign n3052 = ~n2508 & n3051;
  assign n3053 = pi191 & ~n3052;
  assign n3054 = ~n2535 & ~n3053;
  assign po183 = pi150 & ~n3054;
  assign n3056 = pi004 & n2277;
  assign n3057 = pi211 & ~n3056;
  assign n3058 = ~n1584 & ~n3057;
  assign po187 = n1475 | ~n3058;
  assign n3060 = n538 & n1584;
  assign n3061 = pi212 & ~n3056;
  assign po188 = n3060 | n3061;
  assign n3063 = n485 & n2221;
  assign n3064 = pi213 & ~n3056;
  assign po189 = n3063 | n3064;
  assign n3066 = n487 & n2221;
  assign n3067 = pi214 & ~n3056;
  assign po190 = n3066 | n3067;
  assign n3069 = pi215 & ~n3056;
  assign po191 = n1474 | n3069;
  assign n3071 = pi216 & ~n2978;
  assign po192 = n2974 | n3071;
  assign n3073 = ~pi215 & n1474;
  assign n3074 = pi205 & n3073;
  assign n3075 = pi004 & n2307;
  assign n3076 = pi242 & ~n3074;
  assign n3077 = ~n3075 & n3076;
  assign n3078 = pi150 & n3077;
  assign n3079 = ~pi241 & ~po166;
  assign n3080 = ~pi242 & ~n3079;
  assign n3081 = n487 & n3080;
  assign po209 = n3078 | n3081;
  assign n3083 = ~n1860 & ~n2481;
  assign n3084 = ~pi243 & ~n2481;
  assign n3085 = n1860 & n3084;
  assign n3086 = ~n3083 & n3085;
  assign n3087 = n1860 & ~n2481;
  assign n3088 = pi243 & ~n1860;
  assign n3089 = ~n2481 & n3088;
  assign n3090 = ~n3087 & n3089;
  assign po210 = n3086 | n3090;
  assign n3092 = pi243 & ~pi244;
  assign n3093 = ~pi243 & pi244;
  assign n3094 = ~n3092 & ~n3093;
  assign n3095 = ~n2481 & ~n3094;
  assign n3096 = n1860 & n3095;
  assign n3097 = ~n3083 & n3096;
  assign n3098 = pi244 & ~n1860;
  assign n3099 = ~n2481 & n3098;
  assign n3100 = ~n3087 & n3099;
  assign po211 = n3097 | n3100;
  assign n3102 = pi045 & pi046;
  assign n3103 = pi047 & n3102;
  assign n3104 = pi048 & n3103;
  assign n3105 = pi049 & n3104;
  assign n3106 = pi050 & n3105;
  assign n3107 = pi051 & n3106;
  assign n3108 = pi129 & ~n3107;
  assign n3109 = ~pi129 & n3107;
  assign po212 = n3108 | n3109;
  assign n3111 = pi049 & n3103;
  assign n3112 = pi050 & n3111;
  assign n3113 = pi051 & n3112;
  assign n3114 = pi048 & ~n3113;
  assign n3115 = ~pi048 & n3113;
  assign po213 = n3114 | n3115;
  assign n3117 = pi050 & n3103;
  assign n3118 = pi051 & n3117;
  assign n3119 = pi049 & ~n3118;
  assign n3120 = ~pi049 & n3118;
  assign po214 = n3119 | n3120;
  assign n3122 = pi050 & n3102;
  assign n3123 = pi051 & n3122;
  assign n3124 = pi047 & ~n3123;
  assign n3125 = ~pi047 & n3123;
  assign po215 = n3124 | n3125;
  assign n3127 = pi051 & n3102;
  assign n3128 = pi050 & ~n3127;
  assign n3129 = ~pi050 & n3127;
  assign po216 = n3128 | n3129;
  assign n3131 = pi045 & pi051;
  assign n3132 = pi046 & ~n3131;
  assign n3133 = ~pi046 & n3131;
  assign po217 = n3132 | n3133;
  assign n3135 = ~pi045 & pi051;
  assign n3136 = pi045 & ~pi051;
  assign po218 = n3135 | n3136;
  assign n3138 = pi206 & ~n2534;
  assign n3139 = ~pi206 & n2534;
  assign po219 = n3138 | n3139;
  assign n3141 = pi160 & n2531;
  assign n3142 = pi161 & n3141;
  assign n3143 = pi159 & ~n3142;
  assign n3144 = ~pi159 & n3142;
  assign po220 = n3143 | n3144;
  assign n3146 = pi161 & n2531;
  assign n3147 = pi160 & ~n3146;
  assign n3148 = ~pi160 & n3146;
  assign po221 = n3147 | n3148;
  assign n3150 = pi157 & pi161;
  assign n3151 = pi158 & ~n3150;
  assign n3152 = ~pi158 & n3150;
  assign po222 = n3151 | n3152;
  assign n3154 = ~pi157 & pi161;
  assign n3155 = pi157 & ~pi161;
  assign po223 = n3154 | n3155;
  assign po039 = ~pi032;
  assign po050 = ~pi045;
  assign po091 = ~po000;
  assign po112 = ~pi157;
  assign po133 = ~pi021;
  assign po135 = ~pi175;
  assign po151 = ~pi190;
  assign po168 = ~pi205;
  assign po184 = ~pi191;
  assign po185 = ~pi210;
  assign po186 = ~pi039;
endmodule



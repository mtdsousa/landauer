// Benchmark "alu4_cl" written by ABC on Sun Apr 22 21:42:56 2018

module alu4_cl ( 
    pi0, pi1, pi2, pi3, pi4, pi5, pi6, pi7, pi8, pi9,
    po0, po1, po2, po3, po4, po5  );
  input  pi0, pi1, pi2, pi3, pi4, pi5, pi6, pi7, pi8, pi9;
  output po0, po1, po2, po3, po4, po5;
  wire n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
    n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
    n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
    n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
    n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
    n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
    n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
    n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
    n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
    n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148,
    n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
    n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172,
    n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
    n185, n187, n188, n190, n191, n192, n193, n194, n195, n196, n197, n198,
    n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
    n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
    n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234,
    n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
    n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258,
    n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
    n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282,
    n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294,
    n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
    n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
    n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
    n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
    n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
    n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
    n367, n368, n369, n370, n371, n372, n373, n376, n377, n378, n379, n380,
    n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
    n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
    n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n416;
  assign n17 = pi4 & pi5;
  assign n18 = ~pi6 & n17;
  assign n19 = pi0 & pi6;
  assign n20 = ~pi0 & ~pi2;
  assign n21 = pi6 & pi9;
  assign n22 = ~pi7 & ~pi9;
  assign n23 = ~pi6 & n22;
  assign n24 = ~n21 & ~n23;
  assign n25 = ~pi5 & pi6;
  assign n26 = pi5 & pi9;
  assign n27 = pi6 & ~pi7;
  assign n28 = n17 & n27;
  assign n29 = n26 & ~n27;
  assign n30 = ~pi4 & n29;
  assign n31 = pi4 & ~pi9;
  assign n32 = pi7 & n25;
  assign n33 = n31 & n32;
  assign n34 = ~n30 & ~n33;
  assign n35 = ~n28 & n34;
  assign n36 = pi4 & ~pi5;
  assign n37 = pi0 & pi2;
  assign n38 = pi5 & pi7;
  assign n39 = ~pi6 & ~n38;
  assign n40 = ~pi9 & n39;
  assign n41 = pi0 & ~pi2;
  assign n42 = ~pi4 & ~pi5;
  assign n43 = ~pi0 & pi2;
  assign n44 = ~n17 & ~n42;
  assign n45 = pi7 & ~n44;
  assign n46 = ~pi6 & n45;
  assign n47 = pi9 & n46;
  assign n48 = ~pi5 & n27;
  assign n49 = ~pi4 & n48;
  assign n50 = ~n47 & ~n49;
  assign n51 = n37 & ~n50;
  assign n52 = n27 & n43;
  assign n53 = ~n41 & ~n52;
  assign n54 = n26 & ~n53;
  assign n55 = ~pi0 & n40;
  assign n56 = ~n54 & ~n55;
  assign n57 = ~pi4 & ~n56;
  assign n58 = ~n24 & n36;
  assign n59 = ~n20 & n58;
  assign n60 = ~pi2 & ~n35;
  assign n61 = ~n59 & ~n60;
  assign n62 = ~n57 & n61;
  assign n63 = ~n51 & n62;
  assign n64 = ~pi4 & pi5;
  assign n65 = pi6 & n17;
  assign n66 = ~pi6 & ~n63;
  assign n67 = pi6 & n63;
  assign n68 = ~n66 & ~n67;
  assign n69 = ~pi4 & pi7;
  assign n70 = n26 & n69;
  assign n71 = pi9 & n27;
  assign n72 = pi0 & ~n63;
  assign n73 = ~pi0 & n63;
  assign n74 = n70 & ~n73;
  assign n75 = n17 & n72;
  assign n76 = n36 & n37;
  assign n77 = n42 & n63;
  assign n78 = ~n76 & ~n77;
  assign n79 = ~n75 & n78;
  assign n80 = n71 & ~n79;
  assign n81 = ~n74 & ~n80;
  assign n82 = pi0 & ~pi4;
  assign n83 = ~pi6 & n37;
  assign n84 = n70 & n83;
  assign n85 = n36 & n71;
  assign n86 = n81 & n85;
  assign n87 = ~n84 & ~n86;
  assign n88 = n19 & n63;
  assign n89 = pi7 & n88;
  assign n90 = pi0 & ~pi7;
  assign n91 = ~pi6 & n90;
  assign n92 = ~n89 & ~n91;
  assign n93 = ~n17 & ~n92;
  assign n94 = ~pi0 & pi7;
  assign n95 = ~pi7 & n81;
  assign n96 = ~n94 & ~n95;
  assign n97 = n65 & ~n96;
  assign n98 = ~pi0 & ~pi7;
  assign n99 = ~pi4 & n25;
  assign n100 = n98 & n99;
  assign n101 = ~pi6 & pi7;
  assign n102 = n64 & n87;
  assign n103 = n101 & n102;
  assign n104 = ~n100 & ~n103;
  assign n105 = ~n81 & ~n104;
  assign n106 = n17 & n63;
  assign n107 = n81 & ~n87;
  assign n108 = n64 & n107;
  assign n109 = ~n106 & ~n108;
  assign n110 = ~pi6 & ~n109;
  assign n111 = ~pi6 & ~n42;
  assign n112 = ~pi0 & ~n111;
  assign n113 = ~n63 & n112;
  assign n114 = ~n110 & ~n113;
  assign n115 = pi7 & ~n114;
  assign n116 = ~pi6 & n82;
  assign n117 = ~pi5 & n116;
  assign n118 = ~pi7 & n25;
  assign n119 = pi4 & ~n87;
  assign n120 = n118 & n119;
  assign n121 = ~n117 & ~n120;
  assign n122 = n63 & ~n121;
  assign n123 = ~n41 & ~n43;
  assign n124 = pi4 & ~n123;
  assign n125 = ~pi6 & n124;
  assign n126 = n81 & n82;
  assign n127 = ~pi7 & n126;
  assign n128 = ~n125 & ~n127;
  assign n129 = ~pi5 & ~n128;
  assign n130 = n64 & ~n68;
  assign n131 = n25 & ~n63;
  assign n132 = pi4 & n87;
  assign n133 = n131 & n132;
  assign n134 = ~n130 & ~n133;
  assign n135 = ~pi7 & ~n134;
  assign n136 = ~n129 & ~n135;
  assign n137 = ~n122 & n136;
  assign n138 = ~n115 & n137;
  assign n139 = ~n105 & n138;
  assign n140 = ~n97 & n139;
  assign n141 = ~n93 & n140;
  assign n142 = pi9 & ~n141;
  assign n143 = pi4 & ~pi6;
  assign n144 = ~pi4 & pi6;
  assign n145 = ~pi2 & pi6;
  assign n146 = ~pi6 & n63;
  assign n147 = ~n145 & ~n146;
  assign n148 = pi4 & ~n147;
  assign n149 = ~pi7 & n148;
  assign n150 = pi6 & ~n63;
  assign n151 = n43 & n143;
  assign n152 = ~n150 & ~n151;
  assign n153 = ~n82 & ~n144;
  assign n154 = ~n41 & n153;
  assign n155 = n152 & n154;
  assign n156 = pi7 & ~n155;
  assign n157 = ~pi4 & ~n68;
  assign n158 = ~n156 & ~n157;
  assign n159 = ~n149 & n158;
  assign n160 = ~pi5 & ~n159;
  assign n161 = pi5 & n37;
  assign n162 = ~n19 & ~n161;
  assign n163 = pi7 & ~n162;
  assign n164 = ~pi4 & n66;
  assign n165 = pi5 & n69;
  assign n166 = ~n164 & ~n165;
  assign n167 = pi2 & ~n166;
  assign n168 = n20 & n27;
  assign n169 = ~pi4 & n168;
  assign n170 = n37 & n144;
  assign n171 = pi6 & n72;
  assign n172 = pi4 & n171;
  assign n173 = ~n170 & ~n172;
  assign n174 = ~n169 & n173;
  assign n175 = pi5 & ~n174;
  assign n176 = ~n167 & ~n175;
  assign n177 = ~n163 & n176;
  assign n178 = ~n160 & n177;
  assign n179 = ~pi9 & ~n178;
  assign n180 = pi8 & n142;
  assign n181 = ~pi8 & ~n142;
  assign n182 = ~pi7 & n18;
  assign n183 = ~n181 & ~n182;
  assign n184 = ~n180 & n183;
  assign n185 = pi9 & ~n184;
  assign po0 = n179 | n185;
  assign n187 = ~pi5 & n143;
  assign n188 = n37 & n187;
  assign po3 = pi1 & pi3;
  assign n190 = ~pi5 & po3;
  assign n191 = n27 & n190;
  assign n192 = ~pi1 & ~pi3;
  assign n193 = ~pi6 & po3;
  assign n194 = pi1 & ~pi3;
  assign n195 = ~pi1 & pi3;
  assign n196 = ~n31 & n191;
  assign n197 = pi4 & n26;
  assign n198 = pi9 & n42;
  assign n199 = ~n197 & ~n198;
  assign n200 = n193 & ~n199;
  assign n201 = ~pi4 & pi9;
  assign n202 = ~pi5 & n19;
  assign n203 = n201 & n202;
  assign n204 = ~n200 & ~n203;
  assign n205 = pi7 & ~n204;
  assign n206 = n43 & po3;
  assign n207 = pi5 & n195;
  assign n208 = ~n43 & n207;
  assign n209 = ~n206 & ~n208;
  assign n210 = n27 & ~n209;
  assign n211 = n43 & n192;
  assign n212 = ~n43 & n194;
  assign n213 = ~n211 & ~n212;
  assign n214 = pi5 & ~n213;
  assign n215 = ~n210 & ~n214;
  assign n216 = pi9 & ~n215;
  assign n217 = ~pi1 & n40;
  assign n218 = ~n216 & ~n217;
  assign n219 = ~pi4 & ~n218;
  assign n220 = n36 & ~n192;
  assign n221 = ~n24 & n220;
  assign n222 = ~pi3 & ~n35;
  assign n223 = ~n221 & ~n222;
  assign n224 = ~n219 & n223;
  assign n225 = ~n205 & n224;
  assign n226 = ~n196 & n225;
  assign n227 = n72 & ~n226;
  assign n228 = ~n72 & n226;
  assign n229 = ~n227 & ~n228;
  assign n230 = pi1 & ~pi4;
  assign n231 = pi1 & ~n226;
  assign n232 = ~pi1 & n226;
  assign n233 = n70 & ~n232;
  assign n234 = n17 & n231;
  assign n235 = n42 & n226;
  assign n236 = n36 & po3;
  assign n237 = ~n235 & ~n236;
  assign n238 = ~n234 & n237;
  assign n239 = n71 & ~n238;
  assign n240 = ~n233 & ~n239;
  assign n241 = pi0 & ~n81;
  assign n242 = ~n240 & ~n241;
  assign n243 = n240 & n241;
  assign n244 = ~n242 & ~n243;
  assign n245 = n63 & n226;
  assign n246 = n81 & n240;
  assign n247 = n17 & n246;
  assign n248 = ~n25 & ~n144;
  assign n249 = ~n42 & n248;
  assign n250 = n70 & n193;
  assign n251 = n85 & n240;
  assign n252 = ~n250 & ~n251;
  assign n253 = ~n63 & ~n87;
  assign n254 = ~n81 & ~n87;
  assign n255 = pi7 & n192;
  assign n256 = ~po3 & ~n255;
  assign n257 = n188 & ~n256;
  assign n258 = ~pi5 & ~pi6;
  assign n259 = n230 & n258;
  assign n260 = pi1 & ~n249;
  assign n261 = pi7 & n260;
  assign n262 = ~n259 & ~n261;
  assign n263 = ~n229 & ~n262;
  assign n264 = ~n194 & ~n195;
  assign n265 = ~n37 & ~n264;
  assign n266 = pi3 & ~pi7;
  assign n267 = ~n265 & ~n266;
  assign n268 = n187 & ~n267;
  assign n269 = n64 & ~n226;
  assign n270 = pi1 & ~n17;
  assign n271 = ~n269 & ~n270;
  assign n272 = ~pi6 & ~n271;
  assign n273 = pi6 & n245;
  assign n274 = ~n63 & ~n226;
  assign n275 = ~n273 & ~n274;
  assign n276 = n64 & ~n275;
  assign n277 = ~n252 & n253;
  assign n278 = n252 & ~n253;
  assign n279 = ~n277 & ~n278;
  assign n280 = ~n226 & ~n279;
  assign n281 = n252 & n253;
  assign n282 = ~n252 & ~n253;
  assign n283 = ~n281 & ~n282;
  assign n284 = n226 & ~n283;
  assign n285 = ~n280 & ~n284;
  assign n286 = n36 & ~n285;
  assign n287 = ~pi1 & n42;
  assign n288 = ~n244 & n287;
  assign n289 = ~n81 & ~n240;
  assign n290 = n17 & n289;
  assign n291 = ~n247 & ~n290;
  assign n292 = ~n288 & n291;
  assign n293 = ~n286 & n292;
  assign n294 = pi6 & ~n293;
  assign n295 = ~pi5 & n244;
  assign n296 = n230 & n295;
  assign n297 = ~n294 & ~n296;
  assign n298 = ~n276 & n297;
  assign n299 = ~n272 & n298;
  assign n300 = ~pi7 & ~n299;
  assign n301 = n229 & ~n249;
  assign n302 = ~pi0 & n17;
  assign n303 = pi6 & n302;
  assign n304 = ~n301 & ~n303;
  assign n305 = ~pi1 & ~n304;
  assign n306 = ~n252 & n254;
  assign n307 = n252 & ~n254;
  assign n308 = ~n306 & ~n307;
  assign n309 = ~n240 & ~n308;
  assign n310 = n252 & n254;
  assign n311 = ~n252 & ~n254;
  assign n312 = ~n310 & ~n311;
  assign n313 = n240 & ~n312;
  assign n314 = ~n309 & ~n313;
  assign n315 = n64 & ~n314;
  assign n316 = n17 & n245;
  assign n317 = ~n315 & ~n316;
  assign n318 = ~pi6 & ~n317;
  assign n319 = n66 & ~n226;
  assign n320 = pi1 & n19;
  assign n321 = ~n319 & ~n320;
  assign n322 = n17 & ~n321;
  assign n323 = ~n318 & ~n322;
  assign n324 = ~n305 & n323;
  assign n325 = pi7 & ~n324;
  assign n326 = ~n300 & ~n325;
  assign n327 = ~n268 & n326;
  assign n328 = ~n263 & n327;
  assign n329 = ~n257 & n328;
  assign n330 = pi9 & ~n329;
  assign n331 = ~pi4 & ~pi6;
  assign n332 = ~n226 & n331;
  assign n333 = ~pi8 & n142;
  assign n334 = n330 & ~n333;
  assign n335 = ~n330 & n333;
  assign n336 = ~n182 & ~n335;
  assign n337 = ~n334 & n336;
  assign n338 = pi9 & ~n337;
  assign n339 = ~pi3 & pi6;
  assign n340 = ~pi6 & n226;
  assign n341 = ~n339 & ~n340;
  assign n342 = pi4 & ~n341;
  assign n343 = ~pi7 & n342;
  assign n344 = ~pi7 & ~n226;
  assign n345 = n144 & ~n344;
  assign n346 = pi6 & ~n226;
  assign n347 = ~n194 & ~n346;
  assign n348 = n143 & n195;
  assign n349 = ~n230 & ~n348;
  assign n350 = n347 & n349;
  assign n351 = pi7 & ~n350;
  assign n352 = ~n332 & ~n351;
  assign n353 = ~n345 & n352;
  assign n354 = ~n343 & n353;
  assign n355 = ~pi5 & ~n354;
  assign n356 = pi1 & pi6;
  assign n357 = pi5 & po3;
  assign n358 = ~n356 & ~n357;
  assign n359 = pi7 & ~n358;
  assign n360 = ~n165 & ~n332;
  assign n361 = pi3 & ~n360;
  assign n362 = pi4 & n231;
  assign n363 = pi6 & n362;
  assign n364 = n27 & n192;
  assign n365 = ~pi4 & n364;
  assign n366 = n144 & po3;
  assign n367 = ~n365 & ~n366;
  assign n368 = ~n363 & n367;
  assign n369 = pi5 & ~n368;
  assign n370 = ~n361 & ~n369;
  assign n371 = ~n359 & n370;
  assign n372 = ~n355 & n371;
  assign n373 = ~pi9 & ~n372;
  assign po1 = n338 | n373;
  assign po2 = po3 | n192;
  assign n376 = pi5 & n144;
  assign n377 = ~pi7 & n376;
  assign n378 = ~n18 & ~n377;
  assign n379 = n245 & ~n378;
  assign n380 = ~pi1 & ~n241;
  assign n381 = ~pi4 & ~n380;
  assign n382 = ~n240 & n381;
  assign n383 = n226 & ~n253;
  assign n384 = ~n252 & ~n383;
  assign n385 = ~n226 & n253;
  assign n386 = ~n384 & ~n385;
  assign n387 = pi4 & ~n386;
  assign n388 = n230 & n241;
  assign n389 = ~n387 & ~n388;
  assign n390 = ~n382 & n389;
  assign n391 = n25 & ~n390;
  assign n392 = ~n18 & ~n247;
  assign n393 = ~n391 & n392;
  assign n394 = ~pi7 & ~n393;
  assign n395 = ~n240 & ~n307;
  assign n396 = ~n306 & ~n395;
  assign n397 = ~pi6 & ~n396;
  assign n398 = n64 & n397;
  assign n399 = n72 & ~n232;
  assign n400 = ~n231 & ~n399;
  assign n401 = ~n249 & ~n400;
  assign n402 = n188 & ~n192;
  assign n403 = n187 & po3;
  assign n404 = ~pi0 & ~pi1;
  assign n405 = n65 & n404;
  assign n406 = ~n403 & ~n405;
  assign n407 = ~n402 & n406;
  assign n408 = ~n401 & n407;
  assign n409 = ~n398 & n408;
  assign n410 = pi7 & ~n409;
  assign n411 = n330 & n333;
  assign n412 = ~n410 & ~n411;
  assign n413 = ~n394 & n412;
  assign n414 = ~n379 & n413;
  assign po4 = pi9 & ~n414;
  assign n416 = ~n20 & ~n37;
  assign po5 = po2 & ~n416;
endmodule


